��   ��A��*SYST�EM*��V9.1�060 11/�14/2017 A 	  ����DRYRUN�_T  4 �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L �ESTOP_�DSBLAPOW�_RECOVAO{PR�SAW_� �G %$IN�IT	RESUM�E_TYPEND�IST_DIFF>A $ORN41p� d =R�4&�J_  4 �$(F3IDXX��_ICIg�MIX_BG-<y
_NAMc gMODc_USd~�IFY_TI�� �MKR-�  $LIN�c   "_S�IZc�� �. �X $USE_FLC 3!�:&iF*SIMA7#Q�C#QBn'SCAN��AX�+IN�*I���_COUNrR�O( ��!_TMR�_VA�g# h>�ia �'` ����1�+WAR��$�H�!�#Nf3CH�PE�$,O�!PR�'Ioq6��OoATH-� P $ENA#BL+�0B�T���$$CLA�SS  �����1��5��5�0V�ERS��7  ���6|/ �55���E����@MF�0�1RE��%�1{O��wOİO����#EI2.K �O__1_ C_U_g_y_�_�_�_�_ �_�_�_	oo�O)W�?H9@ ,��\k1v\kkljm��1� 2.I  4%� �o�o'  OA_A%�o �o2D#hzY� �����
��� @���0�c$"+ �kdK�@����RA��XOA�1@fNʏ܏�  ��$�6�H�Z�l�~� ����}lLD_A��_A֟ �����0�B�T�f��x����������4JM
�OA�cC!2�l ���/�A�S�e�w��� ������ѿ������ (�:�L�^�pςϔϦ� �������� ��$�6� H�Z�l�~ߐߢߴ��� ��������2�D�V� h�z���������� ��
��'�@�R�d�v� �������������� #�<N`r�� �����& 1J\n���� ����/"/-? X/j/|/�/�/�/�/�/ �/�/??0?3h�4�0 v�g?@