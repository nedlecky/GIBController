��   �A��*SYST�EM*��V9.1�060 11/�14/2017 A 	  ����PASSNA�ME_T   �0 $+ �$'WORD � ? LEVEL � $TI- OUTT4&F/�� $SE�TUPJPROG�RAMJINST�ALLJY  $CURR_OަUSER�NU�M�STSTOP�_TPCHG �V LOG_P NT��N�  6 C�OUNT_DOW�N�$ENB_�PCMPWD� �$DV_� IN�� $C� CR5E��A RM9� =T9DIAG9(|�LVCHK >FULLM/��YXT�CNTD��MENU�A�UTO+�FG_wDSP�RLS��U�BURYBAqN�!eENC/�  CR�YPTE � �4�$$C�L(   ��A�K!�� T @ V� �IONH(�  ���$D�CS_COD?����O%�  W�z'_� �/�(S  JJ*�� L �&�A�91�"K!	? 
 $R!�� =?$?2?H?V?l?z? �?�?�?�?�?�?�?
O� O.ODO���#SUP
� �*�FOXO�#F�xO�O�O�� � �L�A��_ �� �� V�[_t&��j���D�O`_��W_��t ��V�_cGLUGH �1K) t �)�_�_	oo-o ?oQocouo�o�o�o�o �'�_�o�o!3E Wi{�����o ����/�A�S�e� w������������� ��+�=�O�a�s��� ������͟܏��� '�9�K�]�o������� ��ɯ؟د���#�5� G�Y�k�}�������ſ ׿�����1�C�U� g�yϋϝϯ������ ��	��-�?�Q�c�u� �ߙ߽߫�������� �)�;�M�_�q��� �����������%� 7�I�[�m�������� ��������!3E Wi{����� ��%