��   -�A��*SYST�EM*��V9.1�060 11/�14/2017 A   ����CELL_G�RP_T   �� $'FRA�ME $M�OUNT_LOC�CCF_METH�OD  $C�PY_SRC_I�DX_PLATF?RM_OFSCt�DIM_ $BA{SE{ FSETC���AUX_OR�DER   ��XYZ_MAgP �� ��LENGTH�T�TCH_GP_M�~ a AUTORA�IL_4�$$�CLASS  O�����D���DVERSIO�N  ����8LOO�R G��DD<Z$?���q���M,  1 <DYX< [�����C���i�����iO/a/s/�A/�/�/�/$ ��/�/�/	;�$MN�U>A>"�  	 <i!/Q?�A? ?e?w?�?�?�?�?�? �?�?3OO+OMO{OaM���@���.�A3��@�A-C�U[�B�DT�B<?�O��ObO�O*_�5NU/M  ���a��-WTTOOL�%?\ 
�H����=�~��{�u�A3�K�Q��A��PBH  B1�_5]�S�.���R>6T��  �`�_ ;_'o�_/o]oCoUowo �o�o�o�o�o�o�o 	+Y?a�u�@�I_�TcS[mZ_ 