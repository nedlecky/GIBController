��  	p��A��*SYST�EM*��V9.1�060 11/�14/2017 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ��4�AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�>#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO"  � A�LM�"ENB���&ON�!� MDG�/ 0 $DEBUG1A�"d
�$3AO� ."��!�_IF� P $ENABL@QC#� P dC#U5K�!MA�B �"��
� OG�f d� �APPINFwOEQ/ ��L A ?1R5/� H0f69EQUIP 20�NAM� ��2_�OVR�$VE�RSI� ��Q1C�OUPLE,  w $�!PP_D0OCES0�!�81�!�"PC> [1	 �� $SOFT��T_ID�2TO�TAL_EQ� �$@%@NO(BU SPI_INDE]�=EX�2SCREE�N_�4�2SIG��0�?�;@PK�_FI0	$�THKY�GPAN�E0D � DUMMY1d�D�!�EU4�A Q0RG1R��
 � $TIT1d ��� �Dd��D� �D�@�D5�F6��F7�F8�F9�G0 �GW�A�EW�A�E.W�18W �FLW1VW2�aR�!SBN_CF��! 8� !J� ; 
2f1_CMN�T�$FLAG9S]�CHE"� �� ELLSETU�P � $H�O�0 PR<0%�3cMACRO?bR'EPRHhD0D+<@�bb{jdo0UTO�B U�0� 9DEVIC&�CTI�0�� @�13��`Bce#VA�L�#ISP_UN9I��`_DO�f7�iFR_FZ@K%D1�3�A�c�C_W�A�d�a+zOFF_��0N�DELXxL�F0�a�Acq�b?�adp�C?�1`yA�E1�C#�s�ATBXt���MO� XsE 	� [MXs���qwREV�BIL�w�!XI� �rR 7 � OD5`��$NO�PM@��pQ0
� �/�"@�� +�V��!XX@}D�T p E �RD_E
��q$�FSSB�&$CH�KBD_SE�eAUG� Gj2 "_�HTB��� Vxt:5}�8C� �a_EDu �� � C2�2A`S8p�4%$l ttO$OP\@Bbqn!�_OK��US�1P_C� !��d�U ^S`LACI�!Ra�e���� �aCOMM� �0$Da�w�H@�dp ��O�B�@BIG�ALLOW� �(KD2�2e@VA�Rݕd!PAB �`BL8#@S � ,K�a���`S+p"@M_O�]"���CCG�XpN�! $��_ID��`��$�� B�)AS|� c�CCBDD�!{�I����LPz�84_ �CCSCH�1` OcOL��`�MM��zS�C�s$MEA�P�\t�`Tg`�!��TR1Q�a�CN�����FS3k��!/0_�F��( )��p��U�� �!B ���CFn�T X0GR�0���M�qNFLIx�u�@UIRE�x���!� SWIT=$�(�N'`S�"CF_�LIM� �; I@EEDð!�Դ�PT�cp�PJ�dV��&$E��.�`7`�>�ELBOF� ��2ŷ2�p/0ӲSCPdֲ� F�!;�F_��G� �A0WA'RNM pP����P�س��NST� CO�R-���`FLTR^��TRAT TR�>� $ACC�a���� ��r$ORIأ.&��RTj`_S�Fg�@CHGx@I���Tp�A�I� �T�������� �а�"a���HQDh�Rqu�2�BJ; ��C�ц�3��4��5���6�� ��8��9��!X�O�S <� i�{���3�2�ЯLLEC���rMULTIr
2ʓyA|
26�CHILD���
1��B@T_�R w 4� STY2pbܖ=�)2ܐ�8w�s��� |A06$����`�
��meTO2��E��EXT���?��B�f2G2n0r�ƴ�0����R.'k�B  �u���  �"��/% 9a���ð�cQ�s��A!����A��?�M�� =�  q�}�" L0��� ��zcpAM�$JOBꗰ����/�IG}�# d{�*<��-'����u���Z���_M���b$ t{�FL�j��BNG�AgTBA��w��Ɂ/1�@k�j0W� @3P�`X40�|�%��$���t�at��
2J��_)R��W�C�J�*�J�D/5C���`�� n@#�S�P_v`�5¼ & \0RO�O�6# (�S��O_NOM_�`n#@$jc(N"
�w0U�@P�X� ��'�@�� ��1P%)���RA@@���2�"����
$TF,a"�D3S�T
�pQU�16�%�&�!H�b�W�T1:EI!������A���A���A�#Y�NTP��PDBG�DED�(r�P�U��@����ӂ��AqX=�[uTAI�c�BUF��:�m1�a)c �а~6��PIӄ�(� P�7M�8M�
Ip0FF�7SIMsQS�@�KEELCPAT�����"f2�#(?2'���C�*���p�w`JB{��vaDE�C�JQ��E\���+c ������MPL�G$G� �G��_0<jc��1_FPW%0TCV_�3j`سT�#��V��V��Q��HVJR �V�SEG�FRA��O��N S�TRT°N��ySP!Vs�"-1q4,G�&〙R��~R"ryBc-` +����ŻQ ��F��P�@'`�bd'�i�ASIZ�,�7d�fT!c� ;j_i�QRSINF���@S±@F[�l_P�h%PjPL�80�@�fCRC���CCm��d_P�hQ��RۢINwQ�xD�a�eD����6yCE{��7Uyp��Jv� �xE�V�v��F�q_7UFװN�v[P�A��Tx�+��,݀�S1�,1V'SCA��0A$�|!(�A
�ʰ.`�	��/�MARGh����F�nP6�QD±��PL I���[Z��q����wBR\�/� ����.E�� �HwANC+�$LG���O��1{��0��(�AGRC_� K#�@R��,S8�ME]A��9��0f3�RA@�8�AZV ����%O�FCT h�Z�PV"�S~@�ADIٛO٘Y�� Y��X�˔��c�\�qG����BMP�T�V`Y:#�A��AES�:`�s� ҁI��0  �`I�i��DA15ҜP㦗��wB}UI@MMENU9��2W�TITU�b��%sqQh2Z_Qp��#3 x{0Q�$�C�K�S�NO_HEADE,�Z��ͱ���@�����D4�R�r�c�IRTR�@ ��1OERRL��:�5",�Q��OR�R$��>�x�P� "�UN_O/�>T�$SYS��IDhᵧ�?���EV�#|e�|�BPXWO�`z:�6� $SK�!��2΀��T�TRLn9�7 �qAC�P���S�IND�DJ$�� _%��1a����m�PL�Q�BWA���E��D?1��L1�Sb�o�UMMYi9޲��1?� i0�DB��9�8��1PR�a 
}�X�g��9�9 @��$��$Na�LB��:�l�p:�;+�."�PC9�<J�\��ENEq@TF�=�i�p�t��RECO]RD�>H��C�п 9$L��:$��2s��ۀP��Q�ڱ_D��0ROS5�2SK˰4�R�D�`��k ���PA��|x�RETURN�!sMRVU5Q C]R��EWMrRD@�GNAL��2$L�A {�X!;$P��`<$P��� =��?1pC��J#pDO�P�a����r�֟GO_AW@ ��M�O��:�}�CS�S��STCY ?`t�P��ID��t�2�2'�N��O�n�x �pI�� �@ P $zR�B)b��PI'�PO��I_BYZ���yT�b_�HNDGD�A HO��A��P��DSBLw���h(�J@��_�LSG�aB��I@�0	FB5e�FE��zY(�_��cG�Cy0$DO�A�S�MC�@�# PID�YT�H��W� yb#ELE��D�`p���� D Tq�8૓INKR _5U0 L��HA7�=a&�`$�3�`��}��H�E �C�MDL� 2D� .0 G&tW%Cu�W%tJG#�b�W"�b�� ��A �"� 	|�{ev_�SLAVF�F�RIN�0���3��_�m�GP�P�p�@ ����Ҡ�Ҡ�����1bˠa"��`#IDp�]&b�]&W2�$NT�V�3b"VE�4��S�KI��Q�SiC�'2��R�AJ�v�Ac�8TS�AF� U 4_SV>�EXCLUM�Ѱ���ONL�@E3Y�y����HI_V��U�PPLY��Rbq�H@X's3_M�}q�VRFY_i�zq2M��$IO�@����6�`1�R�4�#O���v5LS,�F���4�tA�2(�hP;�P��$��6A"CN��PF�;E(� CN�gCHD���_�Ц���AF CP�#[DT��B#�2 H���"�TA�P��K�� \����I oD $ӐBAg�C!�`�F_60�LH�C���E`K�J��K�j�s$�BmI ���_SG�p K �qCURX�u�� K�jQ��@�b��nX�>~VANNUNc�DE �S(�iP�Ѱ�����Y�Q�`�Z�V"EF���Ic�L @O�F�RǤ�`OTx������
C�¯�Eޱ EM NI%�M�Ub�urUbA\!sdDAY��LOAD����Nb���5ޱ�EFF_WAXI$N�����H�O�`p�f�Z�_
��QG�O�@�ɰ�`
��cE���c�em�NB���a���A8^��aG�P 0�Q2q`H�2q���DUx����8�CA� �QbD���H��IDLE_PW��-u�q��V��V_-pm� ��DIAG��R߀ /$Vx�SE��T����q��� �zD���R�ҏa�V�7�PSW�ӱ �p�p<��emO��a3OH�eJqPP��IR��B��r� �z���P~��Bw�r  ��x���numQB�`���uRQDWg�M	S�@݅AC�O���LIFEh��S�@���N��r#��Q��r�C�SC;��@��NrY�Yɠ=�FLAqC�QOV�/������SUPPOH�E���i�_��tUR�_XP1����ᾗZ��W���;���&�����"�XZ�_A���Y2�C" �T���uNG��t�"ICTm�S }`q�CACHElf�b�:vUN3�⇰SU7FFI��a h���Ĭb��6�°`DwMSWT�T 8�PKEYIMAG@�TM��<��JRܥ$"8A��a� VIE$�^awU BBGL�$�P~#?�J����@Ƥ�V�@� ST� !H���P���P�N`P�<�`P�EMAIg�x|a��xAFAUL%ұW��O�AX��U�� ��pT���qXO< $���S-pv�pIT�BUFu��~!u�e�N`1�SU	B紐�C}$��f�*�SAV2����p5� 3�.�M�Y0�VP9Đ��%���_��m`�ɣOT
�� [sP�0M0�%�ĽB��AX_�`b�0X�'3f�_G��
 YN_o�_`Y�:rD����n�M�Yri�T@FA�F�`DT��� ^aZ"g0G�a&hS��?я   �Z Y�^a[����xѯ���C_�� K��R�� �Rء�ՠ�x�DSPd�x�P���IM2� ����Ex��pU�ׅ�4���M��IP�#x�2X�Dt���TH4�S��Ҹ`T2���HSD=I��ABSC�$C��pVz���_È����dNV11G��4�$���F��d��:Ќ��(�SC�r����M�ERl4x�FBCM�Pl3w�ET� m\΢FU��DU۰2	��6CCD��R�������`R;A^a]`�Bq�meq��ePSp��Ct���C6R��n��_`^H *��LY ��h@���� �P� �#���A��Ca��@Na���a������7���8I	9�������1�
1
1!
1.
1�;
1H
1U
1b
2Rp
2��
2
2!
U2.
2;
2H
2U
U2b
3p
3��3�
3!
3.
3;
3*H
3U
3b
4p��EXT�q^a_ < }p���F����!�<'���u�FDR�t`TǰV@����z!���REM�pF�/�OVM�Ӡ%Aީ)TROV�)DTl=��*MX�,IN�)8[��*�qIND� -��
8s��$DG@����� >�#�	�D�f�� RIV�@G�/�G�EAR��IO �K�"-�N:Ї8�a���0�����.�Z_MCM\���F��U&P�_`a ,~�
�?� 4Q/��0�?�1E�p�1t�$��	�o"b��ȀP����pRI������ET�UP2_ c �k��TDz�Qq�T��P�1SGME�VBBAC�d TF�VB^ԅ)X�%c��)�IFI[���	������E�PT&����F�LUIT�e �]q���UR���a�@JFр��P�s�`I�$u$!RS�@?x-P�J[�CO����VR�T  `x$SHO8�a�P��ASS���8I�B�J$BG_��Q ��Q�Q!�Q.�`^�CDATA�qf�KFU�11?��T2?�pf!�A4��qg |#0wNAV���!P�QR�� S��G�$�VISIT0��SCF��SE@mPXuV3`O�q�aB�B�Abp^Kf$PO`If��FMR2l%h y"b��r z!lЌf~'�?�?�?�&(���u�"_pQ>�pGIT_�AL��pM>6|c?u=DGCLF\�oDGDYUxLD�1BA45+�8?:�/AM\ �V�i��i T��FS��Ƥj P�+ �rl��$EX_�q�x�q1����f�j�p3�{5�v�G���wek �#0)�SW��OΆDEBUG��TN��%GR\@}�Un��BKU��O1� 7 1�PO�`y��e��8�e�MlPLOYO�ç�SM�`EA���Q0G�_E l� �r@e!TER�MɅm҅oaORI�L�΀n҅t�SM_Y�VB΀o҅�q�P��p҅�qUP�qg� -15rl!P���W�m/`G\�npE�LTO��$US=E] NFIGk�����0D�����S�n$U;FR_�$t�����G��`OTȗ��TqAb�z ړNSTM��PATW�n��PTHJ��E�E>�i�N���ARTZ����pZ������REL2���S�HFTI↑��$�_�XPR(�B�� �$)���pq{ LP��§SHIU�tU�� T�AYLO'��aр�@@cR���Q��T�ERV����Rq�"֗�M�2���@���@RyCA��ASYM8ь����WJ��!0E C �L�RH�Up�M� �$��p�:�P�ޠ,�ᠦORM�M�ck�GR��xdr�Re���������a�PHAPTmI��s�2MAn� ��#�8�QW�Q8�e!sHOlP�tt �ܒX�Ed`b�OC���>�1$OPOd|ь��oS�!ZPSPd� ��R����OU����ePR���ŝ�|<��De$PWRV03IM���R_x��0`�	���UDBJĺL�uA@$H]�!^B�ADDR<&H��AG��[�P�I�l�R6b.�qv H+ S��7a���դ����!S�E�a9c�pHSR�MN�BwH`p�|"�^�R�OL(�P ��K%U�*�RO�P��QND_C��s��Ԟ��ROUP���_�0�R���1��b^� �h�h�!i� h�! h�P�bA4`x2��AVEDc���s����xc:P�P��_D�" ��cR��PRM_z�R
�TTP_s��H�qy (~�OB�J3`IґD$<&L�E���*�pz �� -'L / _1TĮ�|�S����HKRL��HIT���P ��Da��|�[RV_S����G��SS0I$JQ�UERY_FLA���HW\���q{�����INCPU�aO+���P<�D ���C��C� �IwOLN�B| 8+ yR@q@$SL�b�$INPUT_��a$����la �Tn SL��q}y ���3��3���1IO	�F_AS:�r~�@$L�@P��Av�Ja
ҝ��@P�àHY;'I"�A� UOP�u `g<&�"9� @���P������@���
�`M-��A�� р��TA٢W�A lP����ϰ�`	%@��PS&BU�`ID �p��lP0%��/%_��L+"����$��� N|(�`}%�I�RCA_CN�  �� � p�6� CY��EA1�! 4a�,� ���'S�k�<2#��DAY_8 3(NTVA�EG 7�8�+#7SCAӠ7#CL@q8!cQ�8"1`��A�c/�$��%�5N_��C�B� 8"1�@���P���1�K�8 �/!�8�Q 2�# R$�A�A��BFK� LAB�$A�`.*GUNI�AC���ITY��T�
�J* �A� X�@lBP�D>Q* R�@pAD�d��AJ'R�AFL�p�P�`
�Ccs
�U�JRwe� �� F��p��>P���BDl3g$J7B�bJ8Y!7�2R(W7)F	Py8?YQAPHIpp�QS\WD�pJ7�J8�uPL_KE~U@  �Ke �LM�! � <ƃ0XR8 �#WA?TCH_VAPaޠ�RH�FIELDbD�y� �R�u� �`�ޑV
焰�QCTR`6��R�q0LDk�� xb�E�_M�����Dv1�LNT9K���COO��Qf	Nt�PfT�����J}f~�V���L}G"d�� !�)?LG_SIZv�g�`�e�p�f�fFD�hI�h�h���f�hˀ�f �`���c;v�p;v;v��`;vˀ;v<�8�~�_Ґ_CM̓�q�p�z��qF���w�t�`��(�a���a�v�` �v�v�`�wI�x�x`���vˀ�v�`RS�P��  (ۀLN�Q貌s��DEB�qE��PX���U��f��Lo�e�DAU��EA�e dġ����GHe��ABOO~}��� C(�pIT��Մ��$R9E��SCR�p0��)D�� �P�MARGI��� ����HJ���S\�W(��z�JGM��MgNCH�FN�R���K��PRG��UqF������FWD���HL�STP��V`��P@��܀��RS$�H��ћC���o��\���U�ɔ[� �sj�`1��G��7�PO������r���OCU��RGEX.TUI��I p�3 �  q\�?�q�?���UA����u���d��N�	��ANA�dA�VAI@P�e3DeD�CS0�ӻ��ӻ�O���OͷS�#�ظS�?�IGN�`80�cp��`�1ĴDEV^�LL�qÁX#�`i��Pf!T�r$�g�]H3�d�b�A8����P�0� >��U$۠1��2��3��p�@S»��`� ��)�d�녜0%��`��۠�(Q�STy�R��Y��A� �$EP�CP�P��_�r�P��a� L % 7SpL.L�0���-����֔��_ � �Y��Q3�	��
�MCY��� �� CLDP|yDeTRQLINA��F5�#�FLGTcLD��W�c1D�QW� �LDW�A�W�ORG��A[�j�xRESE�RVF��R��] ��� �,`A�[��2�W�SVI�5�B	�����RCLMC&�����8�h �Q�QM�� o��P�c�MA6d	0�3}r��Tԡ�&%E)PTpa��MISC�E� d,b���RQ�B	tPu`�	0�@� ��(���AX�Db�P��	EXCE%S1����M�n��f@��Dd����S}C�� � H�1��_�0��� u:�Kk� \w@/d���B_�PFLIC���B��QUIRE�i�j`�O��f$L��ML��Mj� ���� b.c&����NDw�� ��`�W��h_D�ss�INAUT�s��`Py�NpbSq�Et��MPSTL�Q� �4�0LOC��RI�P@��EX�ANGx�b����ODAQ�Uŝ��&B�@}RMF b�e&&���&���L%�T���SUP����F�X�@IGG� � �,`��SqO4��s����PaP%@Ӕ)C� �(Cг&� ݣ�1|��1��2��X TpM�@}� t MD1DB) 6��*4=�'7H�Q�*4DIA.A+3�@W�N�*4���*5D��)�O�C�P� H CU�`Vh0Y����OA�_x�Q� ������#z�b���`�8P�>/�P�0P��8KEu��P�s-$qB�p�6��ND2?�S+A2_TX��XЛ@��WBQ�� LOģ��P�FmD�B�lFZ���2�F�C4R�R2�E�` &�}A��A� d$OCALI��TuG��:�G2��RIN�q�Cw<$R�@SW0D��SQ�ABC%(D_�J=@��@1_J3:2V
,R1SP�P}0�@P,TS]3R]�1��
�@�UJQ�U����OZ�IMQ�a�CS�KPD��T�p8c�TJ��a�Q�\�U�U�U�W��_AZ�Q$aE�L?��R?�OCMP0�b�4�k�RT��Oc�E1��PmE��1��qh`�jZ}dSMG�>�0_�JG��SCyL) �SPH_�a��p�c4��@�@R'TERP�C��@9_���sGRAA�8��a�tDI:ab��I-N�`ACT��2$udB��1
#q��_N�A��1uLr
vLHua�Vyvj@DH) d@�A���$V�@x�c`�$�`���������4���R�3�@�H �$BEL5`�e�a_ACCEL����xQ��IRCi_pi��NT4ў �$PS�p(�L  �6�=�$p�!����"A�yo��o�3>�� ,_���r��������CS��p_MGS�$DDÁr��FW�0�s߅��r�ԈDE��PPABmNF�RO�`EE�� ��-�5��Q��{�q �q~>�$USE_�@J{�P� C��{�Y���p� ��YN��A �����PA1��M��1̱���OL_���INC�4������ܗ�Q.��ENC�`L�!�2�6��r��3�IN(�I�>�#�0�dNTVEx���C?�23_U�Q���Q�LOWL�`��l05��q�DF�� ���`����C<p8�MOS���0�����`�PERCH  ��OA@�b Ч�ۣ �!t�_��!JgBbw�}�$�SA>�0�Lz��S���W9�l t�o���T3RK�e%�AY�C*� q��>������Ufu�5�MOM�2��q ��0�����G��q�̳³@DU�P��S_�BCKLSH_C >�1ţ�A@���3P���Zʤ��UCLAL�M5��������CH�K5��S��RTY@� C#��՞�1_;�N��_UM����C��pÁ�a��8�LMTOP�_L��=c�Q1�E �6�(��+�1�+�dP0��9�w��PC��!H��ǅ��C4�SD\��ՇCN_�BND�L��Q�SF�q�Vw������a��>���CAT��SHA#�BՄ �����~E?�~Ir`fĀPA��ڒ_P��ɳ_�PЦ�Ġ�Q�����JG% ? ��_��OG���bTORQUi�gU���������a�-�_W����{a@�qL��sK��sK�IS�Ia�I�sF >�RX���Q̀VC�p0��y��1��; ���Q���JRK�����0D�B�`M�3�0Mv_sDL�qJ�GRVR�`K�sK�s,H_�C8*r�y
COS�W`�LN �����p �	�`�	}��
���'1Z� ��,MY�%�$A�FTHET=0z�NK23�spl�c� CBuCB�cC�@AS�!�}���s�uSB�s��'GTS�Q8�CVQ���ug��g��$DU��S�!"�B���1&ĸQ��Q�"����NE
�T^�K��aix�pdAh�%�'x���LPH�o"I�o"S ���#��#�o"�3(�*�pV�(V�(�p��,V�*V�+V�+V�;V;V;V-9H��(�&�2�-O��8�+H��+H;H;H;H*-9O�,O�(O^I�.UO�*O�+O�+O;UO;O;OFo"���I��D�'SPB?ALANCE�T���LE�H_hSP�)q�IR�IR�PFULCMXtR\WtR��6z1�QaUTO_<����T1T2�Y�r2N�� �A��Tdqٱ�vPT E��s��T`�O�:`�<�INSEG ���REV�V��2�gDIF��[y1�@g6r1���OB6a|��U�2�A���4L�CHWAR�|�A�B���$MEC�H�5���a��AX���PZ��f�'�r�P�� 
�b*��q�RO�BĠCR>�u�� ��DO_DA�T�q� < ����rc���� BE�q$ON5�Xx_�x����qD��� �/� %�T"�*����T7a��L����C�K����CT1  #%�s(��pNĠ�PLsĠRG����b�u�bX�u,p��MP��E�"? $IR�p���C�b�MAI1 hԑ��(�_qp&��C`!���R@ COD�KsFU��FLAG��ID_c�j�#`	�~)PG_SUFF}�� ����#`��F�rDO�w`�uO��GRqr�s���s���b����b˅�,t  �2�:pHj`_FIvAq9�ORDUq�    MMY�36^�����p$�ZDTq�(qxp/u��4 *BaL_N�Aaq�px��uDEF�_I��x��v���uS	T�Q�uP%a�p�u���uΕ�vISX ��Dq�g �t��s��!�"=�4��q�ΒD�P*=�KsD
�O+PCrLOCKE�ᢃ��0�w	�����UM��x� ������Ε������� ������ޔ��e��� 	����`�῅x����� ���N���{pPh`���p�m �pW��������TEs��0t� �n�ULO�MB_����0�V�IS� ITY�Ar��Oq�FRI�S��i`SI��YAR��pǾp�3���$W�W��< � 9_Y�ɁEASBqsùS��� �Gh��o h �pTEk`�)�7n�COEFF�_O�q%�Ěqp`G$Z�|�Si�k�PvP/pBp �$����W�A�wqGRX  � � $��RMrX�pTMr�&���rX��@�VsER4`Th��g���  �RLL�ʄ�⬡SVB����$��������{ �SETU��wq�4p� � l��+� 6�ID�� �b��W���}��pW�s�T���;�Ԃ*��qP��O�6�F k`EB�R)�3���uq�SK_,P�� �P:pT1_USER�Q���`���QVEL-���`���r�qIQ�7 �MT{q�C���  ��pH`O�bNORE�S^r���OPWO� �,��SY�SBU�0!�SOP(�t� �T#�U"�C`1P���I�PA����XK�b!�OP��U5�=�ha?r5�}�IM�AG���Px�;�IMW��IN< q��?RGOVRDQ09���|�P~��pg >�hC����bL}�BT%">��PMC_EY�(�)�N�@M5�>�1�94�  ���SL�gP� ��`OV�SL�VS}�DEX@3�ܐ`L eq��_�� x���x��>��C�`z��U����?��~� @� Q � �eOr�RIZ��!P�>���EaE�� �H��`|�ATUS>��$TRCY ��DXUB*�bK���-�4�7Y�� D :qz�cU�0�V$���^���XE\�հ������ ��[U1P)����PX���w+�3-�	�P�G���$SU�BJ�e��JJMPWAIT��b%WLOW�bF�qMY��aRCVF6��p�b�e!RE� Fa�qC�� RL�b�p�'IG�NR_PLDB�TB|�P��aBW�V��$��Ump�%IG�a��p�Q�TNLNl�&2RT��NO�yN�pZPEED�>iHADOW|��c��ERVEhV4w�4!��SP�P � L:p�`��v0b�4�UNI��0!R���LYN��PTr<P��~� 0� @��~��p0p9P �NePgKET�2 �BU��PIP�"~Ἕ�ARSIZ[�%��ۑ�<Ò~"ORMA�T�P�$g�BbEM2�d@D�3UX����PLo��� $��r�SWI�`�b���WO�a�e�P�LV�AL_ ���@�0A-�BʰC�-�D�� �,��J3�D�H� T��PD�CK  �!�CO_�J3�PH�CSBaE��.��O�M	���|�!  � �Ep?PAYLOA�CkT�_1rZ2rS�@J3AR��X~U�V�S�_RTIA4�Y5�Y6-�MOM-��S�S��S�S�S{pBy AD��Sf�Sf�SPUB��pR�T9e�S9e�R���E{��� L$�PIV1mS��wUX�j�uWZ�j���j�kI�c�PnQ3��f!�f#!$RO
R�#/r�:3HIG�C:3z% s4-vs4z%� � -vcs�<x�!Ky�!z%SAM�P��1�y-w�sz%M'OV_.����q g�3����t �v��P�y�P��R|��T�uf� fr�u�/�f��s5�Q��,�z"7�w�N�w���GAMM#�S^�^!7GETrFI�3h`4\S��
��IB��2�Ir0C�)�h�Ad���EP����'�LW�T�K�6�@x�'���v0�AC�%GCHK���^#I_�pB���d�kY e����S��f���C� �$�H �1��I��RCH�_D��2� �$4�L�E���m�WX5���0MSWFL�$Mn�PSCR(75�� �t2�\@¥�g��P�y`թ�0��0�ASVna7�P��UR����׏�SAV'���:�C�NO[PCD�\T :��k_�asY�isY �`�����`/R�eԸ�SDO�1A�o��uת �'x�7v!�cx8�4����qD�bdMz�� �йBYL�c�q��ЏЊ��Ƿ ��	������q�𨠷!N�M_Wi����=`���l�M� ��CL�ȱQ�$1�a0�"
���{����$���$W��WANG��Q��3TH�:T H�ATH��D� 4����(�C��p�X�0OBSo��Z��
�� M�� ���OM�uV|���p����Ŀ�PCON`��U�bc[Q_��� | Q�:��Y���S���S�:��Z����Z�A� P��	�x������P�x�P0A�PM� Q}U�p � 8� �QCOU���QT�H� HO��?�HY�SG@ES�q>�UE�*�0�	@O8$�  b�@P� �UN]ʶ��@Or�� �P����%��2ROOGRAp��2�O���ITA0��l��INFOna� ГA������E�OI���� (�SLE�Q�'u' ����OyS��7$� 4� �ENABvҫ PTIONV4�b�j4�[GCFd��JX� o������R�����OS_E9Dg �� �W��ЩK�qL#�E%�N9UAUTV�COPY�qp/!�b�M�N9=��PWRUTj� @N� ;OU�B$G��� �R�@� � � � ��k�T!?USR_TSP3�{TP�KLNA�t�CL��%#T9P
&y	DBG�����9&q8'�1@L�D��]� ��s ��� ASK��4����M�PA9�yP�3�!PRG_� "�!��v�%U@�*K/  ��I\Ѭ$CH�@�(��$ <�_OVzCT� �Z�2MJ�PTICT��}O��STATU;C�I�0f9AP�@h7M�O_WA� r083X �3�0�#���������CR���4?�94�1C6��:R5 6�5/G/�Y/k$2s%�� ,&� HE�b0A�����m`aEg1 1� �WKT(�� <� Nj�TRIE�)"SE)�NC�� 	WE`EQǂ�< r�,�A���. �@�B�G�CLU�2PRIp�B�@�#�WRKz o� �W�SV���,�)VS��t$�5E�XECf9�1�B �jV#�2�@OOF0O �	We �܄&ETELE: 2�{ �GADJna�� h��X� MI�U���f��fWhP�h{�f6s�P83EX_T_CYCv�j�'RGN�0b�x����LGO����NYQ_F�0��W�����a� s��LA}�aa����(�0��J���IF1Y��
'�b_G}g3�e~�Ma@�rU�qo�:�LASTqT�hd��Qd� �`nFEASIq8��rˠ ��Mr8C�v3B��� �B���b.aB��r��r�AB)!�E��2�VAq�vBASO��v��Ο�UPDǁO��$�q �RMS_T�R�so�`����SP�J�:q �VjbM��:��	�U� ���� ��q�
�p�?�'�n���p
����e�DOU��[��2hdPR]��P۞.GRID��)#B�ARS�&zr�ROsTO�!�� y�D�!!!1`�TO��.a� ��L)�w�R�%B�k�_�SA�)`�X�DIX�T_ �Pz���]���P��l �������6��7��8�x�j�F�C�P�w�$VALU�s-�qt�o��@F`�� !mQ���*�!*�b AN,��q�!Z1U�TOTA�$s�p�|�PW�cI߁��R�EGEN������X����Z5�F�%�TR�sr��_S0�󧤠��sVa�T��S�qE�&s�D�T�X�V_H �DA%��V�GS_Y���ҧfS=�{AR%�2� ��I1 E;���X�6u_@��1�^Q�����ip���&ͫ��SLG��
d� {q�f�2)�d0$pS��7tDEw�1U{q~���TE���P�� !̡B;�J�7C�cIL_�M�d��V�r���T!Q%�#���C�氂5V��C��P_���p���M��V1��V1���2��2��3��3
��4��4�ʻ�Pu�`��]y��!v�IN�ٟVIB11�Ŧ�2���2��2��3��3
��4��4�؜Я�������B�D $�MC_FH��`A	2 ��nl�M��0�1=�1⸃ �ก�E�Vh�$KEEP_HNADD*��!l��pv�CCOM��!���+�|p��O �k�s)� ��g1�c��REb0��#q�B�������U
$e��HPWD  l��SB�"1�COLL�AB!�?��m��b�q2�0O�����T�=�R@$FLp��q�$SYN#�z�M��C�����UP_WDLY ��p�LA��$qqBY��A�DX��4�Q�SKIPk�� �,�D�OR��T�Ѣ����RR����O�p� �p�Q	]	�Q	 l!	ǐ
Ԑ
�
t�
9-a�RA)��� X��S�f�MB�LIC�#� �0U��&Sw�0�A��q^W�SWIT�� �_� AMGV�� ��XQ\u$U�W�J0�/��:�NGRLT��O�s��,�.�8�1*�T_Jl! �}5R_WEIGH��#J4CHq`VOqR�V3�LOOe���r�qTJC�(�EcA0�e��OB�pY5?
$C�J2� ��-�ɲEX�pT�c!ITW�!� h�!ұ�h�f`RDCQ�n��� �PR3�TOR�@����R�af*�q�<g s�RGEA좠pm#��FLG�p0~�Ts�SPC+"�5 >j�2TH2NQ�|!y@� ����POS11��� �l]���/�&P�A�T���1U�53IN�4,20s�,2U��oHOMEW2 
222�??1?C?�U?g? �� 332���?�?�?�?�?�? � 24B�OO+OP=OOOaOy75B�O��O�O�O�O�O C
�$6B�__%_7_�I_[_ �%7B��~_�_�_�_�_�_ M 28B��_oo�1oCoUoy5S0����  2� 3��� ��3��@G��ɰ0� rr�sIOg�-y�I�`opsCPOWE��� �`��:!��$$C��=S� ���zq� ��  opC�SIܡ�xw�p����$AAVM_�WRK 2 zu� 0  �5�q��x���} �|	 !��5�� {p�#�`�G�e������ ���0ˏݏ儩pBS�0S!� 1�y� <��*�<�N�`� r���������̟ޟ� ��&�8�J�\�n��� ������ȯگ���� "�4�F�X�j�|����� ��Ŀֿ�����0� B�T�f�xϊϜϮ��� ��������,�>���}C��AXLMTqvA���  dS��IN\�n�R�PRE�� E��Ў���C�_U�O  �z� ��C߶�ID ?yzu�� � ��&�8�a�\�n��8�����SET�ؾq��� ���UPDAT�����  �pI�OCNV_� � �j�P3�1�
����8� 1�{P $���K�������{p?��aж������� ��"4FXj| ������� 0BTfx�� �����//,/ >/P/b/t/�/�/�/�/ �/�/�/??(?:?L? ^?p?�?�?�?�?�?�? �? OO$O6OHOZOlO ~O�O�O�O�O�O�O�O _ _2_D_V_h_z_�_ �_�_�_�_�_�_
oo .o@oRodovo�o�o�o �o�o�o�o*< N`r����� ����&�8�J�\� n���������ȏڏ� ���"�4�F�X�j�|� ������ğ֟���� �0�B�T�f�x������S�LARMRECOV �eю��o�LMDG ��������_I�F �f�d$�SRVO-053� Disturb�ance exc�ess(G:1 �A:3) ,1 �d Root H�ub f#0, �ut#9�����d�����ÿտ��, �
�� 5����8�CHECK_SL�OT C�LINE� 0C�AUTO ABORTEDC�C�JOIN~�rτ���NGTOL  ���	 A  � ����S�PPIN�FO �� ��� ��$�6�e�  
�8�f��Uߏ�y� �ߝ߯���������C����o��� ������������#��5�G���PPLIC�ATION ?�(����Handli�ngToola� �
V9.10P�/05��R�
1�4203P©�42�95609��16�57��������7�DF1��R�C�No�neR�FRA�R� ��_�_A�CTIVE��  �x��  uV�M�OD ���rCHGAPONL���� OUPLEDw 1&�� � ��lCUREoQ 1	&�  p�$$	u�|� ��Wi{�����/���$���$H�p��(*HTTHKY</�/*/0/�/ �/�/�/�/�/??n? 8?J?\?z?�?�?�?�? �?�?�?�?OjO4OFO XOvO|O�O�O�O�O�O �O�O_f_0_B_T_r_ x_�_�_�_�_�_�_�_ obo,o>oPonoto�o �o�o�o�o�o�o^ (:Ljp��� ���� �Z�$�6� H�f�l�~�������Ə ؏���V� �2�D�b� h�z�������ԟ� ��R��.�@�^�d�v� ��������Я���N���*�<�Z�`�r�6T�O����DO_C�LEAN�s��N�M  �� �$G�Y�k�}Ϗ�*D?SPDRYR �rHI� #�@4���� �1�C�U�g�yߋߝ�p������oMAXf� ങ�s����X�������uPLUGGp� ���PRC��B!�%�����K��OP����SEGF� K����!�3������1�C�{��LAP����U#�������� ����'9K]|o�TOTAL�|<�USENU���� Ƹ�s�6R�GDISPMMCʷ��C���@@$���O��������_STRING �1
�
��M� Sq

F_�ITEM1P  nql~���� ���/ /2/D/V/�h/z/�/�/�/�/�I/O SIGN�ALJTry�out Mode�QInp0SimulatedU�Out<O�VERR�� = �100TIn �cycl5UP�rog Abor�3U�$Stat�usS	Hear�tbeatOM?H Faul�7�3Aler�9�/�?�? �?�?OO/OAOSOeO ܳLܱ^hO �O�O�O�O�O_"_4_ F_X_j_|_�_�_�_�_p�_�_�_|OWOR�� L2a�OoZolo~o�o �o�o�o�o�o�o  2DVhz���~POJ�1�pJk� ���/�A�S�e�w� ��������я������+�=�O��rDEV �~z��g�����şן �����1�C�U�g� y���������ӯ���PALT�M�Jo ��F�X�j�|������� Ŀֿ�����0�B��T�f�xϊ��GRI ��L��6��������  �2�D�V�h�zߌߞ� ����������
��.��Ϩ R�Mf���@�� ������������� 0�B�T�f�x�������x����T�PREG"�  ~���2DVhz �������
�.@Rdv�-��$ARG_2`D �?	������  w	$�&	[��]���'��SB�N_CONFIG�� �12!C�II_SAVE � �$+!""�T�CELLSETU�P �%  ?OME_IO�-�,%MOV_Ho �/�/REPi��/�UTOBACKZ!��("UD1;:\�� �/@'/   q0��#8��C139��18/02/2�8 06:58:34������?�?�?�?<���?O(O :OLO^OpO���O�O �O�O�O�O�O�O_._ @_R_d_v_�__�_�_ �_�_�_o�_*o<oNo�`oro�o�ou��  �1_�#_\ATB�CKCTL.TM�P G.DG L��p�/�o�o�/I�NI!�V5&�#MESSAG: DqE!�� #VtODE_ADt =&%.!zuO|����#PAUS�q!��� , 	������w,		���<�&�8� r�\�������̏�����ڏ��&��t�pTSK�  �}#?)� UgPDT}pBwd����vXWZD_ENqBBt*��STAAu�����XIS U�NT 2�+!�D � 	 9�u�!���� ��{�?����&�����  �  ��  �u��E0�  ��R�d�&���E0�, v�� _x �p ��C���g����گݔMETh�2�I�F# P��EE�bE!X@ET��VC�X�D����E�Tj��;�?2;k�/<�p��;܇s;�.�<.����SCRDCFG �1�1 	�87D ǯ������ ѿ���?��U4:�� F�X�j�|ώϠ���� +�������0�Bߩ��ϥ�!GR吇����Ӹ`NA� �	��$}�_ED@p1�k�� 
 �%{-�`EDT-n���*	SCAN_S#LOAp�\�]'$� Q-�#������?x�&�ߝ�  ����A2��+����b�QF5 B��'�n������!3_������R�?耈���:�L���p���4 +�+	���<�T� �<��5�g D�� ���z��6�3/W���W/��F/���7 �/��/#/��/#?j/|/?�/��8[?���?������?�?6?H?�?�l?��9'O�?tO�?� ��PO�OOO�O8O��CR���/?_Q_ =_��_�O�Ot__����N�O_DEL��~�GE_UNUSE���|�IGALLOW� 1��   �(*SYST�EM*��	$S?ERV_GR�Ҷ��?`�pREGHe$8jc��?`NUMmj�c��mPMU�P���LAY�����PMPAL�?CYC10�^�nq�`�nsULS'�`�o`f�b�qJcL~TtBOXORIqe�CUR_Ap�mPoMCNV�fAp�10�n�pT4DL�I��:\i	*PR�OGRAGdP�G_MI�n�	�AQL�u� �	�B4��?n$FLUI_RESU�gm�wo��\�_��̏ޏ�� ��&�8�J�\�n��� ������ȟڟ���� "�4�F�X�j�|��������į֯���]X��L�AL_OUT �.ki��WD_A�BOR�`oa�IT�R_RTN  �D���d�NONS�TO�Џ� hC�CG_CONFIG ��������� �°E_RIgA_I`��(����°FCFG �������1�_�LIMVb2��= �`� 	fߗϢ�B<bҴ��e�@��`�PAN�GP 1];������)�;���CH`\�n�+C1r�9r�@rЯ��C��CVr�]r�d
r�lr�sV�����߫C[��mr�vr��rЄrЈ� C�jrБ�Ж�G?����HE�Pɳm��G_�P�p1��  �U��`�r��������
�HKPAUSf^q1��(� �b� �	������}��A��U5������ (+���N� ��:�x�^��������� ������>$b4t°O5�;�Q�~�LLECT_5�ao�X�JǱEN�pp��v���NDE��o�c�R1�234567890!�BYaK�1�C'
 H#��C)l� Y\k}�4���/ ��/f/1/C/U/�/ y/�/�/�/�/�/�/>? 	??-?�?Q?c?u?�?��?�?�?O1��i��� ��IOG !
�����`�O�O�O�ObGTR��#2"FM-�}I
�?�N�̰#qMZT��_�MORi�$�� �>��A����U ���Y�_�_�_�_�_�[�dR��j�%r],�?$��>c��KHd����P�'�U� ߔo�o�o��
�o�o R�ޱ�ƾȍ�r"��o��� �Q!\XP�DB� )L�Dc?pmidbg5�LO�s:��>wqp||��v  ��>1z��}���la��}�>�mgR���v��~f���Z��>@ud1:�A��ZZqDEF (�R|C),�cQ�b?uf.txtL��|\M�Xp_MCkS*L��TC�����jT+Ν�|T�K�A���Cf�Bf��C�CC�3k�B�fC��\C!H�C��ǭ�ʅ�D����Di�oD����E+�\D�w�IEv��F�F����F���F���HG?��F�)�Gc�ʾ�>Cc������g-FL��R���EU`XZ�����D���)x�+���о���3D��fE�̅��EX�EQ��EJP F�E��F� G��n�^F E�� �FB� H,- Ge��H3YE�;?����33���#v  n�r�Q#5ٛ��R��AAa��=L��<#�SU��.п���RSMOFST &k��v��P_T1�D�E .fo��XQ����;�ɲ���?���<��M��TESTe�,k�)�R�/����KC4���j� ����Cz$��"��Ъ"�C�@�E�^Sa:d�
��I%0��?VӸ�1r]I��:�RT_e�PR/OG k%����|��j@NUSER�����KEY_TB�L  ��~`�u�	�
�� !�"#$%&'()�*+,-./*:�;<=>?@AB�Ce�GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~�������������������������������������������������������������������������������͓���������������������������������耇��������������������6A��LCK���������STAT+���_A�UTO_DO���_�IND�N��1RK�j�\�T2�����STO:��� TR�L��LET�����_SCREEN� rZkc�sc � U��MMENU 12a{ <�ܵ�}�e \������� �-c:Lr ������/�  /&/_/6/H/�/l/~/ �/�/�/�/?�/�/I?  ?2??V?h?�?�?�? �?�?�?�?3O
OOBO {OROdO�O�O�O�O�O �O�O/___e_<_N_ �_r_�_�_�_�_�_o �_oOo&o8o^o�ono �o�o�o�o�o�o�K"4��<_M�ANUAL��ZCD\�3����������߿�?|(�t�s��4�� B�~���$DBCO���RIG5�b�_E7RRL��5Λa������� G��NUMLI��������U�DBPXW�ORK 16Λ����0�B�T�f���D�BTB_�� 7�v��ڑ��E�D�B_AWAYO�^GCP ��=x���_AL��N���K��Y��������i� �18�� , 

�����9�v���K_M��I�Ȝ@�����ONTIMM�������
����MOTNEND����RECORDw 1>�� �~���G�O�F�4��� ɒr�������?���׿ F���j��1�C�ڿ� y�违���������� ��ߊ�?߮�c�u߇� ��߽�,���P��� )�;��_��߃��ߧ� ������L��p���� I�[�m�������� 6�����!��E0 >{�����2� �h�ASe� t�
�.��/ ��=/�a/��ru �/�//�/�/S/?w/�� ��/B?T?�/��TOLERENCǔsB��ՐL��G��CSS_CNST_CY 2?�����	`?���?�?�?�? OO0OBOXOfOxO�O �O�O�O�O�O�O__��4DEVICE ;2@�; ��j_ _�_�_�_�_�_�_�_�o!o��3HNDG�D A�;�Cz�4j��1LS 2BT]3o�o�o�o�o�o��o5o�2PARAM C��v�r�e~teRBT 2E���8d�<q_���Ck�v0  � !~������3�B��w!uB�O  ��w���~܀�y���g�,��|A�!sC�0l�(���K�pZ�A��!u�H!vc�}!v�x� ��̏�����&�8��J���n���͟�2�){�Df`C�0��� 	 AZff�Aa��A��0
:������ff!z��MC�Car�!��*��D�,��Bo���Bj��B3J���ffB���C%CL��"�4�F�(���;m� ڠ��!} �s����ꯥ�ӯ��� 	��h�?�Q���u��� ������Ͽ���R� )�;�M�_�qσ��ϧ� ���ߓ�0�B�-�f� Qߊ�u߮ߙ����߿� ����,���b�9�K� ��o��������� ����L�#�5�G���k� }������� ������ H��lW���� �������) ?Q�u��� ����/R/)/;/ �/_/q/�/�/�/�/? �/�/<??%?7?�?� �?�?�?�?�?O�?&O OJO%S?e?�OM?{O �O�O�O�O_�O�OF_ _/_A_S_e_w_�_�_ �_�_�_�_�_oo+o xoOoao�o�o;O�o�o �o,PbM� aO�o�o����� ��L�#�5���Y�k� �������� �׏�6� ��l�C�U�g����� ���e� ��D�/� h�S���w���¯�˟ ݟ
���@��)�;� M�_�q���������˿ ݿ���%�r�I�[� ��ϑϣϵ�����&� ��J�5�G߀�kߤߏ� �߳�����ٯ���� �/�|�S�e���� �������0���f� =�O�a�s��������� ����b�߆ q�������(&
�$DCSS�_SLAVE �F���W��@_4D � WlCFG �GWa;d�MC:\JL�%04d.CSV�64�  �?A� �CH�z@ ��/7/=  ��FT!d/R)Q!X�N���#C.?�@ E)�RC_O_UT HW�"�;_C_FSI �?W �+�??1?Z?U? g?y?�?�?�?�?�?�? �?	O2O-O?OQOzOuO �O�O�O�O�O�O
__ _)_R_M___q_�_�_ �_�_�_�_�_o*o%o 7oIoromoo�o�o�o �o�o�o!JE Wi������ ��"��/�A�j�e� w���������я���� ��B�=�O�a����� ����ҟ͟ߟ��� '�9�b�]�o������� ��ɯ�����:�5� G�Y���}�����ʿſ ׿����1�Z�U� g�yϢϝϯ������� ��	�2�-�?�Q�z�u� �ߙ��߽�����
�� �)�R�M�_�q��� ����������*�%� 7�I�r�m�������� ������!JE Wi������ ��"/Aje w������� //B/=/O/a/�/�/ �/�/�/�/�/�/?? '?9?b?]?o?�?�?�? �?�?�?�?�?O:O5O GOYO�O}O�O�O�O�O �O�O___1_Z_U_ g_y_�_�_�_�_�_�_ �_	o2o-o?oQozouo �o�o�o�o�o�o
 )RM_q�� ������*�%� 7�I�r�m�������� Ǐُ����!�J�E� W�i���������ڟ՟ ���"��/�A�j�e� w���������ѯ���� ��B�=�O�a����� ����ҿͿ߿����'�9�b�]�o��$D�CS_C_FSO ?������ P u�oϸ������� � )�$�6�H�q�l�~ߐ� �ߴ��������� � I�D�V�h����� ��������!��.�@� i�d�v����������� ����A<N` �������� &8a\n� �������/ 9/4/F/X/�/|/�/�/ �/�/�/�/???0? Y?T?f?x?�?�?�?�?��?�?�?��C_RPI����OUO~OyO $O��HO�O�O�O�O��SL6O@�O
_S_|_ w_�_�_�_�_�_�_o oo+oToOoaoso�o �o�o�o�o�o�o, '9Kto��� ������#�L� G�Y�k���������܏ ׏���$��1�C�l� g�y���������ӟ�� ��	��D�?�Q�c��� ������ԯϯ��� �"_�OF_(�q����� �����ݿ��*�%� 7�I�r�m�ϑϺϵ� ��������!�J�E� W�iߒߍߟ߱����� ����"��/�A�j�e� w����������� ��B�=�O�a����� ������������ '9b]o��� �����:5��LPRE_CHKg J�KLA L��< ��Q�E���E 	 <���Y��/-/ /Q/c/=/O/�/�/�/ �/�/�/??�/?M? _?9?�?�?o?�?�?� �?OO�?7OIO#OUO OYOkO�O�O�O�O�O �O	_3___i_{_U_ �_�_�_�_�_�?�?o /o�_;oeo?oQo�o�o �o�o�o�o�o�o Oa;��q�� �����9�K�o 3�����m���ɏ��� ��ُ�5�G�!�k�}� W������������՟ �1��U�g�]�O��� ��I�ӯ寿����� �Q�c�=�����s��� Ͽ�������;�M� '�Yσ�y�������e� �������7�I�#�m� �Yߋߵߏߡ����� ��!�3��?�i�C�U� ������������ /�	�S�e�?�����u� ����������= O);��q�� �����9K� o�[����� ��#/5//A/k/E/ W/�/�/�/�/�/�/�/ ?'U?g??s?�? w?�?�?�?�?	OO�? 'OQO+O=O�O�OsO�O �O�O�O_�O�O;_M_ '_q_�_=?k_�_�_�_ �_o�_%o7oo#omo oYo�o�o�o�o�o�o �o!3WiC� ��_������ �)�S�-�?�����u� ��я��ݏ���=� O�)�s���_������ ������9��%� o���[�������ï� ǯٯ#�5��Y�k�E� w���{���׿�ÿ� �ٟ�U�g�Aϋϝ� w����ϭϿ�	���� ?�Q�+�u߇�a�s߽� �ߩ������)�;�1� #�q�������� ������%�7��[�m� G�y���}��������� !��-WM�_� �9���� �AS-_�cu ����/�/=/ /)/s/�/_/�/�/u �/�/?�/'?9??]? o?I?[?�?�?�?�?�? �?O#O�?OYOkOEO �O�O{O�O�O�/�O_ _�OC_U_/_a_�_e_ w_�_�_�_�_	o�_o ?oo+ouo�oao�o�o �o�o�o�O�O);�o GqK]���� ���%���[�m� G�����}���ُ��ŏ �!���E�W�?��� ��y�ß՟������ ��A�S�-�w���c��� ����������+�=� �a�s�i�[�����U� ߿�˿��'���]� o�Iϓϥ�ϱ��ϵ� ���#���G�Y�3�e� �߅�������q���� ����C�U�/�y��e� ��������	���-� ?��K�u�O�a����� ����������); _qK����� ��%�I[5 G��}���� /�E/W/�{/�/ g/�/�/�/�/�/?�/ /?A??M?w?Q?c?�? �?�?�?�?�?O+O!/ 3/aOsOOO�O�O�O �O�O�O_'__3_]_ 7_I_�_�__�_�_�_��_o�_�_GoYo����$DCS_SG�N KIE�`��3"w620�-NOV-18 ?14:35 ;c�`�8-FEB�a07�:53�`�`�b� L\>��aMF3MaO-�a�b�i�`�aq߀��7[bC��w9��o  qcVERS�ION }jV4.2.0|�EFLOGIC �1LIE�  	:`�fN@�ayN@p~CrPROG_ENB  �d�Xs�`�sULSE�  vu�uCr_�ACCLIM�v���s��sWR�STJNT�w�a�mdEMO�|�a�q�Br�INIT �MPzEJ�OPT?_SL ?	IF'��
 	R57Y5�c{�74��6���7��56t��1��2���bxϏ=w^�TO C j��o$�>vV5��DEX�wd�b�`�<�PATH A�}jA\ YST�EM VOLUM�E INFORM�ATp\*���sH�CP_CLNTI�D ?!vXs �bx�eڟrIAG_GRP 2RIE� �6qQ@D�  �D�� D  �B�  B�6�3ff�j%�B�6�Q���kM��6�y�g����B�N�C�-Bz��Bp6��e`�imp�2m7 7890?123456̡ ��Q@�  Ao��mAj1Ad�A]�
AW�|�AP�AJ�-AC/A;��A4>�頸a@��  A�`A��A,)�U�A�6�6��`;B4�l �ej���a
�uƨAp�ffAj�yAe�K�A_�AYAS��MC��AF��A@ � EJ!�3�E�EJY�ANm��@�X�ȑ�@��y����Ŀ�ֿ����;d��5?@~ff@x�1'@q��@k�C�@d�D@]?��@Vv�,�>��P�b�t���s��l���@e@^���@W\)@O���@H��?2�7K�@.V��������� ���S@M�&�G2�A��@<�1@5��@/�l�@(Ĝ@!���\D�V�h�z� ��n�]oB�AN1�w�� �]���������� ����O�a�?�����!���NC����¡�-Ѽ��@�>��R ?�33?Y�����@�7'Ŭz(6) 4�F4���L@�@�p��P�
=@�O@�Q�`�m@=��Ah�Ф���J�=� c<��]>�*�H>V>�3�>���@�?<���<� ����l֐�?� ��C�  <(��U�b 4L�3a3��� �iA@�b?H���:��Hn� GH���P���x/"/��?�7D!�>�(�>��P!=����@���G�l/G�@����՝%�m����н @����@�`@Q�?LT�����Ũ�I�F�ܦ�e?4��' �p61A?�&��]4g?F��C�  C���CC'o? <�?�? 5e���  94L�6o���4C��18!�6p��8!�?�0�����A�D
�J�`6u㡫?,O(�?PO9lHxH�� I;8j�V��8C3��=H�@O�O<O�O�O	_�O�-_�DICT_C�ONFIG S��)��de�gwu�STBF_TTS�w
�y�Sp�s�a�Vq`MAU��p�rMSW_C5F\PT�  A�z�OCVIEW�PU�]K����AoSo eowo�o�omR/o�o�o �o�o�oBTf x��+���� ��,��P�b�t��� ����9�Ώ����� (���L�^�p������� ��G�ܟ� ��$�6� şZ�l�~�������D\KRC�SV%�R!P� ���!��E�4�i�X�����TSBL_FA?ULT Wߪh>��GPMSK�W���PPTDIAG �X`Y�QoS��UD1: 6�78901234A5�nR�nW��P*_ S�e�wωϛϭϿ��� ������+�=�O�a� s�6�u�
Bϻ�>JVTRECP��
��)��A�>�P� b�t��������� ����(�:�L�^����ߩߦ�gUMP_?OPTION�P��F��TR�R�S�����PME�U��Y_T�EMP  Èϓ3B�pP5 �A2 UNI�P�U5��VYN_BRK �YoMREDITCOR����_�пENT 1Zߩ�  ,&
CH�ECK_SLOT� RAME����&
SCAN_L�ABEL�f�&�UPDATE_B�OXF�FICND mP%	���P
SAFE�Z ��&-BCKEDT- ���&S� 7�$�QUICK �P$!//DE�MO +/e+&MAINR/�/�BG }/�/�GENER�/�/	�&VIZPIX� G 1�/�,L?IGHTIN?�/{N�EST12?�
TOOLY1__?5TOY0� ^?�.�S' �2�?	Z��?O��EMGDI_STAHdQ5mQm � NC7C1[�[� �d�OrO�N
�Nd���O�O�O_!_ 3_E_W_i_{_�_�_�_ �_�_�_�_oo/oAo So��jo|o�o�o�i�A �o�o�o�o
.@ Rdv����� ����*�<��jco m�������oǏُ� ���!�3�E�W�i�{� ������ß՟���� �/�A�[�e�w����� ����ѯ�����+� =�O�a�s��������� Ϳ߿���'�9�S� A�oρϓϭ������� �����#�5�G�Y�k� }ߏߡ߳��������� ��1�K�]�g�y�� A����������	�� -�?�Q�c�u������� ��������)C� U�_q����� ��%7I[ m������ �/!/3/MW/i/{/ �/��/�/�/�/�/? ?/?A?S?e?w?�?�? �?�?�?�?�?OO+O E/OOaOsO�O�/�O�O �O�O�O__'_9_K_ ]_o_�_�_�_�_�_�_ �_�_o#o=O/oYoko }o�O�O�o�o�o�o�o 1CUgy� ������	�� 5oGoQ�c�u����o�� ��Ϗ����)�;� M�_�q���������˟ ݟ�����?�I�[� m��������ǯٯ� ���!�3�E�W�i�{� ������ÿտ���� �7�A�S�e�wϑ��� �Ͽ���������+� =�O�a�s߅ߗߩ߻� ��������/��K� ]�o��������� �����#�5�G�Y�k� }��������������� '�9�CUg�� ������	 -?Qcu��� ����/1;/ M/_/q/��/�/�/�/ �/�/??%?7?I?[? m??�?�?�?�?�?�? �?O)/3OEOWOiO�/ �O�O�O�O�O�O�O_ _/_A_S_e_w_�_�_ �_�_�_�_�_o!O+o =oOoao{Omo�o�o�o �o�o�o'9K ]o������ ��o�5�G�Y�so �o������ŏ׏��� ��1�C�U�g�y��� ������ӟ����#� -�?�Q�c�}������� ��ϯ����)�;� M�_�q���������˿ ݿ�i��%�7�I�[� u�ϑϣϵ������� ���!�3�E�W�i�{� �ߟ߱���������� �/�A�S�m�w��� �����������+� =�O�a�s��������� ���������'9K e�[������ ��#5GYk }������ /1/C/�oy/�/ �/�/�/�/�/�/	?? -???Q?c?u?�?�?�? �?�?�?�/O)O;O MOg/qO�O�O�O�O�O �O�O__%_7_I_[_ m__�_�_�_�_�_�_ Oo!o3oEo_Oio{o �o�o�o�o�o�o�o /ASew�� �����_��+� =�WoI�s��������� ͏ߏ���'�9�K� ]�o���������ɟ۟ ���#�5�O�a�k� }�������ůׯ��� ��1�C�U�g�y��� ������ӿ���	�� -�?�Y�c�uχϙϫ� ����������)�;� M�_�q߃ߕߧ߹��� E�����%�7�Q�[� m����������� ���!�3�E�W�i�{� �������������� /I�Sew�� �����+ =Oas���� ����//'/A7/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?Y?k?�}?�?�?�?�?� ��$ENETMOD�E 1\B%��  ��A�BGK�0�RROR_PRO/G %�:%�aO�nI<ETABLE  �;L/�O�O�O��G<BSEV_NU�M 
B  ��AP<A_AU�TO_ENB  q(EC9D_NOQ� ]�;A R�  *�YP�YP�YP�YPP+XPr_�_<�_2TFLTR_0V�HIS�C�@+[_�ALM 1^�;� ��Y\�+ �_2oDoVohozo�o�_�_�B8P  �;�WQB�j�0TCP_�VER !�:!�YO�o$EXTLO�G_REQ�V�)Y#sSIZ,tSkTKIyGU� r�TOL  �D�z�R�A t_BWD�`�p�V�q#Bv�sDI�q _B%��sD��{S�TEP���0�pO�P_DOk�1FA�CTORY_TU�N�Wd3�DR_G�RP 1`�9�Qd� 	�o��@{���*v���R�HB ��2 ���� �e: ������{�Џ�˄@�_�BO��AT�6���Q!�"���G��� @>������A�@��[�@��A�.dP`���!@F�nA�(A��&@�'�A9��\P8������n�XY�8�?/���@h�A9��?y�?�h��@�њ
 F�5U&��v�Gx��џ	bE�ҟ�D�a�L����B� � ��A����33�33^�UUU�ʪ@��۠j�%G>u�.�>*��<�����E�� F�@ ��&��J���NJk�I�'PKHu��IP�sF!��֞�  j��9��<9�8�96C'6<�,5����g� *�� 8�����} i�7W���tKF�EATURE �aB%�p"A�Handling�Tool 	���English� Diction�ary�4D S�t��ard	��A�nalog I/�O@�I�gle S�hift\�uto� Softwar�e Update���matic B�ackupɯ�g�round Ed�it��Came�raW�F[�Cnr�RndIm����o�mmon cal�ib UI���n����Monito�r&�tr�Rel�iabp��DHC�P�]�ata A�cquis5�^�iagnos��T�x��ocument �VieweA�`�u�al Check Safety!�~�hanced!�4���s��Fr����xt. DIO �1�fi��&�end.��Err@�L��B�J�sA�rR�1� �p��FCTN Me�nu��v\Ӕ�TPw In��fac����G��p Mas_k Exc��g#��HT��Proxy� Sv����igh�-Spe��Ski�����5�mmun�ic��ons �u�r����s�X���connect 2W��ncr��struH#�U�~�e����J����KAREL C�md. L��ua����Run-Ti�"�Env����el� +��s��S/W��License�����X�Book(System)�MACROs,�?/Offsew�:aH5���q�? MR:��6Ҭ�MechSt�op��tn��:iS�s˪x��T���i�odq�witch��~��._�Op�tm~��fil���}gM�:ult�i-T�����PC�M fun���o������Regi�/ r;��ri��F���U�Num S�el�� � Ad�ju+��!!s�2-t�atu�J/���R�DM Robot> �scove)��%em� 5�n7ǆ%�"Servo5�� �?SNPX b��x�;SN��Cli���.t�Libr(�?��Q �0�&o t���ssag��` 0��R��`/I��f5�MILIB�?i2P� Firm��y>PΡ�Acc����TPsTXm�g4elnR �?j1�Nz=orq}uq�imula?�4��*Fu� Pa��y>���Z�&��ev.�f5��ri��OU�SB port ��iPL�a�жEn?except�Ы ���E��VC�r6�-�V��R�?,U4;&[S 0SC�5^_�SUI�Web Pla&�^�!M��T�������x�ZDT Appl4���F�_g�Grid�!pla�ymv0�� gRR.�7�Zf��3_=-10�iA/1r�]�DV�-k�Path C�trîk��eJ�l�arm Caus�e/� ed*ȉ�S��W@rityAv/oidM�l�7�#Gu=�0rP��)�es9�t�c��ycp������@��a�CS �./�c�Ҏx���W�j��therNet�1����q@�1�EDA��xScal�AЖ�RAn@ �Y�v�te  �APMC/�A�Pk��}O:x�����NRTL�?��On�e Hel؊I�C�������Katr;�x 8r��mHap����64MB DRA9M��T�FRO]��Ŝ|��ellW��sh����ȗc/ŕ��YppFڜtyp�s"D���r��rzt��(.xۖus�s��mai��;�ݑ �"T�q��T1��W�OAdp.խ�s����C�}
�L̀ar��!9���:R7�9ayx�d��OPT ��*� !cY0l��&��r w�kپ*5Nd�.
 ��Ouest�%�"S�p�du[��� SWI�MEST f@�4�295609ud� vbM�D�Vσ�zόϹ� ���������
��I� @�R��v߈ߵ߬߾� �������E�<�N� {�r��������� ���A�8�J�w�n� �������������� =4Fsj|� �����9 0Bofx��� ����/5/,/>/ k/b/t/�/�/�/�/�/ �/�/?1?(?:?g?^? p?�?�?�?�?�?�?�?  O-O$O6OcOZOlO�O �O�O�O�O�O�O�O)_  _2___V_h_�_�_�_ �_�_�_�_�_%oo.o [oRodo�o�o�o�o�o �o�o�o!*WN `������� ���&�S�J�\��� ���������ڏ�� �"�O�F�X���|��� ����ߟ֟���� K�B�T���x������� ۯү����G�>� P�}�t�������׿ο ����C�:�L�y� pςϔϦ�������	�  ��?�6�H�u�l�~� �ߢ����������� ;�2�D�q�h�z��� ���������
�7�.� @�m�d�v��������� ������3*<i `r������ �/&8e\n �������� +/"/4/a/X/j/|/�/ �/�/�/�/�/�/'?? 0?]?T?f?x?�?�?�? �?�?�?�?#OO,OYO PObOtO�O�O�O�O�O �O�O__(_U_L_^_ p_�_�_�_�_�_�_�_ oo$oQoHoZolo~o �o�o�o�o�o�o  MDVhz�� �����
��I� @�R�d�v�������ُ Џ����E�<�N� `�r�������՟̟ޟ ���A�8�J�\�n� ������ѯȯگ��� �=�4�F�X�j����� ��ͿĿֿ����9� 0�B�T�fϓϊϜ��� ���������5�,�>� P�bߏ߆ߘ��߼��� �����1�(�:�L�^� �������������  �-�$�6�H�Z���~� ��������������)  2DV�z�� �����%. @Rv���� ���!//*/</N/ {/r/�/�/�/�/�/�/ �/??&?8?J?w?n?��?�?�?�?�?�2 � H552��3�121ER78�H50EJ614�EATUP)F54�5)H6EVCAM�ECRIdGUIFv)G28eFNREF�52XFR63GS{CHEDOCV�FwCSUF869)G�04FEIOC�G4�FR69XFESE�TAGWGJ7WGMA{SKEPRXY}H]7FOCOX3AHhF!P(H3TVJ6'H�53�FH�XLCH^<VOPLGAG0lV�MHCR=VS�WMkCS@H0$W554F�MDSWg_WOP�_WMPR`V�@�X0n(FPCM|FR0[g�!P4F�P�W51LG5u1�h0LFPRSW�69TVFRDdFR�MCNF93(FS�NBA�G�WSHLEB�fMw�@h2(F�HTC@FTMIL�H�FTPA�FTPTXAvEL�f�P�Gq8G@FJ95�F�TUT`W95TVU�EC<VUFRdFV�CC�xO�VVIPNLvCSCpv�@IEwWEB@FHTT@F�R6�H�xCG/�I�G�IPGSU�R�CLvDG_WH77�4FR8g��LFR6m6��51 W53�g[68��66lX2lX�6�h6�FR7kWRc82�y��'H76(F���TVR58��x5�4P�66؈GNV�DVR79 W84ֈFD0�F��RT�S�fCLIDhKGC�MS�F��@FSTY:Lw6gCTO@F�@��FJNNTVORSn�VR68D�53�544wPMDi�W�h�@4FOPIl���WPRQFL�wSJ��SVS�FGene D�8����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{����������� ����/ASe w������� +=Oas� ������// '/9/K/]/o/�/�/�/ �/�/�/�/�/?#?5? G?Y?k?}?�?�?�?�? �?�?�?OO1OCOUO gOyO�O�O�O�O�O�O �O	__-_?_Q_c_u_ �_�_�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o% 7I[m��� �����!�3�E� W�i�{�������ÏՏ �����/�A�S�e� w���������џ��� ��+�=�O�a�s��� ������ͯ߯��� '�9�K�]�o��������ɿۿ�  ?H552���21	�R78�5�0	�J614	�AwTUP9�5459̽6	�VCAM	�C�RI��UIF9�2�8��NRE�52�x�R63�SCH�	�DOCV��CS]U�8699�0HʯEIOC��4�R{69x�ESETY��w�J7w�MASK^	�PRXY��7	�OCOy�3Y�ʅ��8�3��J67�53�(�H�LCH��O�PLGY�0��MH�CR��Sg�MCS�X�0��55H�MD�SW����OP��M�PR�����08�PCM��R0'���H�lu��51h�51h��0h�PRSx�69���FRD��RMC�N	�938�SNByA���SHLB���M����28�HT=CX�TMIL�(��TPAH�TPTXFY
EL��u�(�8'��%��J95��TU�T��95��UEC��UFR��VCC�(O��VIPh
C�SC�
�I	�WE�BX�HTTX�R6l���CG�IGwoIPGS�RCh
�DG��H77H�Rq8��% h�R668+�51X�53X�68V+66��2��6h��6��R7��R82�8,7�768�% ��gR58�,�54;s66x,�NVDxڷR79X�84��Du0W;F�<RTS���CLI�g�CMS�H��0X�STYh6���CTOX��H�J�NN��ORS��R�68;53�+54HPM�x����H��OPI��0(KPR�Q�L7SfLSV=S��Gene	�� O_a_s_�_�_�_�_�_ �_�_oo'o9oKo]o oo�o�o�o�o�o�o�o �o#5GYk} �������� �1�C�U�g�y����� ����ӏ���	��-� ?�Q�c�u��������� ϟ����)�;�M� _�q���������˯ݯ ���%�7�I�[�m� �������ǿٿ��� �!�3�E�W�i�{ύ� �ϱ����������� /�A�S�e�w߉ߛ߭� ����������+�=� O�a�s������� ������'�9�K�]� o��������������� ��#5GYk} ������� 1CUgy�� �����	//-/ ?/Q/c/u/�/�/�/�/ �/�/�/??)?;?M? _?q?�?�?�?�?�?�? �?OO%O7OIO[OmO O�O�O�O�O�O�O�O _!_3_E_W_i_{_�_ �_�_�_�_�_�_oo /oAoSoeowo�o�o�o �o�o�o�o+= Oas����� ����'�9�K�]� o���������ɏۏ� ���#�5�G�Y�k�}� ������şן���� �1�C�U�g�y����� ����ӯ���	��-� ?�Q�c�u����������Ͽ��ST�D�LANG �� �2�D�V�h�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r����� ��������&�8�J� \�n������������� ����"4FXj�|
RBT�OPTN������ );M_q���DPNĿ�� �//+/=/O/a/s/��/�/�/�/�/�+ted ��??'?9? K?]?o?�?�?�?�?�? �?�?�?O#O5OGOYO kO}O�O�O�O�O�O�O �O__1_C_U_g_y_ �_�_�_�_�_�_�_	o o-o?oQocouo�o�o �o�o�o�o�o) ;M_q���� �����%�7�I� [�m��������Ǐُ ����!�3�E�W�i� {�������ß՟��� ��/�A�S�e�w��� ������ѯ����� +�=�O�a�s������� ��Ϳ߿���'�9� K�]�oρϓϥϷ��� �������#�5�G�Y� k�}ߏߡ߳������� ����1�C�U�g�y� ������������	� �-�?�Q�c�u����� ����������) ;M_q���� ���%7I [m����� ��/!/3/E/W/i/ {/�/�/�/�/�/�/�/@??/?A?S?e>�k?��?�?�?�?�?�:9�9�5�$FEAT�_ADD ?	����A@  	�8%O7OIO [OmOO�O�O�O�O�O �O�O_!_3_E_W_i_ {_�_�_�_�_�_�_�_ oo/oAoSoeowo�o �o�o�o�o�o�o +=Oas��� ������'�9� K�]�o���������ɏ ۏ����#�5�G�Y� k�}�������şן� ����1�C�U�g�y� ��������ӯ���	� �-�?�Q�c�u����� ����Ͽ����)� ;�M�_�qσϕϧϹ� ��������%�7�I� [�m�ߑߣߵ����� �����!�3�E�W�i� {������������ ��/�A�S�e�w��� ������������DDEMO aI?   �8N DV�z���� ���I@R v������ �//E/</N/{/r/ �/�/�/�/�/�/�/
? ?A?8?J?w?n?�?�? �?�?�?�?�?OO=O 4OFOsOjO|O�O�O�O �O�O�O__9_0_B_ o_f_x_�_�_�_�_�_ �_�_o5o,o>okobo to�o�o�o�o�o�o�o 1(:g^p� ������ �-� $�6�c�Z�l������� ϏƏ؏���)� �2� _�V�h�������˟ ԟ���%��.�[�R� d�������ǯ��Я� ��!��*�W�N�`��� ����ÿ��̿��� �&�S�J�\ωπϒ� �϶���������"� O�F�X߅�|ߎ߻߲� ���������K�B� T��x�������� �����G�>�P�}� t������������� C:Lyp� �����	  ?6Hul~�� ���/�/;/2/ D/q/h/z/�/�/�/�/ �/?�/
?7?.?@?m? d?v?�?�?�?�?�?�? �?O3O*O<OiO`OrO �O�O�O�O�O�O�O_ /_&_8_e_\_n_�_�_ �_�_�_�_�_�_+o"o 4oaoXojo�o�o�o�o �o�o�o�o'0] Tf������ ��#��,�Y�P�b� �������������� ��(�U�L�^����� �������ܟ��� $�Q�H�Z���~����� ���د��� �M� D�V���z�������ݿ Կ��
��I�@�R� �vψϢϬ������� ���E�<�N�{�r� �ߞߨ��������� �A�8�J�w�n��� ������������=� 4�F�s�j�|������� ������90B ofx����� ��5,>kb t������� /1/(/:/g/^/p/�/ �/�/�/�/�/�/ ?-? $?6?c?Z?l?�?�?�? �?�?�?�?�?)O O2O _OVOhO�O�O�O�O�O �O�O�O%__._[_R_ d_~_�_�_�_�_�_�_ �_!oo*oWoNo`ozo �o�o�o�o�o�o�o &SJ\v�� �������"� O�F�X�r�|������� ߏ֏����K�B� T�n�x�������۟ҟ ����G�>�P�j� t�������ׯί�� ��C�:�L�f�p��� ����ӿʿܿ	� �� ?�6�H�b�lϙϐϢ� ����������;�2� D�^�hߕߌߞ����� �����
�7�.�@�Z� d����������� ���3�*�<�V�`��� �������������� /&8R\��� ������+" 4NX�|��� ����'//0/J/ T/�/x/�/�/�/�/�/ �/�/#??,?F?P?}? t?�?�?�?�?�?�?�? OO(OBOLOyOpO�O �O�O�O�O�O�O__ $_>_H_u_l_~_�_�_ �_�_�_�_oo o:o Doqohozo�o�o�o�o �o�o
6@m dv���������2�   )�H�Z�l�~������� Ə؏���� �2�D� V�h�z�������ԟ ���
��.�@�R�d� v���������Я��� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t� �������������� (:L^p�� ����� $ 6HZl~��� ����/ /2/D/ V/h/z/�/�/�/�/�/ �/�/
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o FoXojo|o�o�o�o�o �o�o�o0BT fx������ ���,�>�P�b�t� ��������Ώ���� �(�:�L�^�p����� ����ʟܟ� ��$� 6�H�Z�l�~������� Ưد���� �2�D� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬϾ������� ��*�<�N�`�r߄� �ߨߺ��������� &�8�J�\�n���� �����������"�4� F�X�j�|����������������0	  1+L^p �������  $6HZl~� ������/ / 2/D/V/h/z/�/�/�/ �/�/�/�/
??.?@? R?d?v?�?�?�?�?�? �?�?OO*O<ONO`O rO�O�O�O�O�O�O�O __&_8_J_\_n_�_ �_�_�_�_�_�_�_o "o4oFoXojo|o�o�o �o�o�o�o�o0 BTfx���� �����,�>�P� b�t���������Ώ�� ���(�:�L�^�p� ��������ʟܟ� � �$�6�H�Z�l�~��� ����Ưد���� � 2�D�V�h�z������� ¿Կ���
��.�@� R�d�vψϚϬϾ��� ������*�<�N�`� r߄ߖߨߺ������� ��&�8�J�\�n�� ������������� "�4�F�X�j�|����� ����������0 BTfx���� ���,>P bt������ �//(/:/L/^/p/ �/�/�/�/�/�/�/ ? ?$?6?H?Z?l?~?�? �?�?�?�?�?�?O O 2ODOVOhOzO�O�O�O �O�O�O�O
__._@_ R_d_v_�_�_�_�_�_ �_�_oo*o<oNo`o ro�o�o�o�o�o�o�o &8J\n� �������� "�4�F�X�j�|����� ��ď֏�����0� B�T�f�x��������� ҟ�����,�>�P� b�t���������ί� ���(�:�L�^�p� ��������ʿܿ� � �$�6�H�Z�l�~ϐ� �ϴ���������� � 2�D�V�h�zߌߞ߰� ��������
��.�@� R�d�v������� ������*�<�N�`� r���������������P&6: - Pbt����� ��(:L^ p�������  //$/6/H/Z/l/~/ �/�/�/�/�/�/�/?  ?2?D?V?h?z?�?�? �?�?�?�?�?
OO.O @OROdOvO�O�O�O�O �O�O�O__*_<_N_ `_r_�_�_�_�_�_�_ �_oo&o8oJo\ono �o�o�o�o�o�o�o�o "4FXj|� �������� 0�B�T�f�x������� ��ҏ�����,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ����  �2�D�V�h�zόϞ� ����������
��.� @�R�d�v߈ߚ߬߾� ��������*�<�N� `�r��������� ����&�8�J�\�n� ���������������� "4FXj|� ������ 0BTfx��� ����//,/>/ P/b/t/�/�/�/�/�/ �/�/??(?:?L?^? p?�?�?�?�?�?�?�?  OO$O6OHOZOlO~O �O�O�O�O�O�O�O_  _2_D_V_h_z_�_�_ �_�_�_�_�_
oo.o @oRodovo�o�o�o�o �o�o�o*<N `r����������&�8��$F�EAT_DEMO�IN  =���h��>�P�IND�EX]�l��P�I�LECOMP �b������k�K���SETU�P2 c��~���  N Ӂ���_AP2BCK� 1d��  #�)9���%��:�>���(�e�;�����  ���D��z���� 3�E�ԟi�������.� ïR���������A� ЯN�w����*���ѿ `������+Ϻ�O�޿ sυ�ϩ�8���\��� ߒ�'߶�K�]��ρ� ߥ߷�F���j���� ��5���Y���f��� ��B�����x����1� C���g������,��� P���t�����?�� cu�(��^ ��)�M�q  ~�6�Z�/ �%/�I/[/�// �/�/D/�/h/�/�/
?�3?���P� 2>��*.VR:?�?� *�?�?�#�?�?��%n0PC�?O� OFR6:�?4N�?XO�;T|�|O�OEyO�L_�IO�O�&*.Fq?_�!	C�O<\q�O`_�KSTMk_ �_B"@�_�]O_�_�KH�_o�Wo�_�_io�JGIFso�o�U��oFoXo�o�JJPG �o!�U�o�oq�:#JS{�� 7s��O%
JavaS�cript��oC�S�(��V�� %�Cascadi�ng Style SheetsT��� 
ARGNAMOE.DT���,�P�\��U��qǄ؏��>ǀDISP*Ώ����P�[��M�\��
�TPEINS.X3ML��7�:\��]����Custom Toolbar����PASSWOR�DR��.FRS:�\#�� %Pa�ssword Configd��/�� <����?���+�=� ̯a�𯅿��&���J� ߿n���Ϥ�9�ȿ2� o�����"Ϸ���X��� |��#߲�G���k��� ߡ�0���T߾��ߊ� ��C�U���y��� ��>���b�����-� ��Q���J������:� ����p���);�� _���$�H� l��7�[m �� ��V�z /��E/�i/�b/ �/./�/R/�/�/�/? �/A?S?�/w??�?*? <?�?`?�?�?�?+O�? OO�?sO�OO�O8O�O �OnO_�O'_�O�O]_ �O�__z_�_F_�_j_ �_o�_5o�_Yoko�_ �oo�oBoTo�oxo �oC�og�o�� ,�P����� ?���u����(��� Ϗ^�󏂏�)���M� ܏q������6�˟Z� l����%����[�� ������D�ٯh��� ���3�¯W������ ���@����v�Ϛ� /�A�пe����ϛ�*π��N���rτ������$FILE_DG�BCK 1d������� < �)
S�UMMARY.DyG#���MD:W������Diag� Summary��ߥ�
CONSLOG��p߂������Console� log��	T�PACCN�v�%�^���TP A�ccountin�=��FR6:I�PKDMP.ZI	P����
�� ��շ��Exceptio�n$���*.DT�S�|���FR:\�g���/�FR DT Files������MEMCHECCK���߆�+/��Memory D�ata,��'?�)	FTP���61�mme?nt TBD�`�o �)ETHERNET�������3��Ethe�rnet 3�fi�guraC��ĚDCSVRF���ܵ<%z v�erify al�l�c�y�uDIFF���:/= �%�diff�</���zCHG011//*/�/�R/�/�?<})2�/�/�/ C?N/�/�/�"39? ?2?�? Y?�?}6�VTRNDIAG.LS�?�?�?KOz>A Ope[� Log ��no�stic`н��)VDEVBD�A��(O:O�O�V�isnADevic9euO�KIMGB�ЪO�OQ_T3�DImsag�O�KUP�@�ES�O,_FRS�:\�_����Upd�ates Lis�t�_��?PFLEXEVEN)0_B_�[o�a UIF� Ev�r@\og r���)
PSRB?WLD.CM�o����R�o�_0�PS_ROBOWEL�
��Iq9Do]�8KNet/I�P�0a�odŎuSMp�L�8��q/Email܆_��l!rSHADOW���i��<Shadow? Chang��a��L!rRCME�RRa�F�X��<���CFG Err�or�@t��� �o��SGL�IB�̏ޏs�>6� St\|A�+�on)_�ZD�p͟\��8ZDq@�ad�� �j��NO�TIП�w�:Notific\ �a�h��ί�� �����(���L�ۯp� �����5�ʿܿk� � ��$�6�ſZ��~�� �ϴ�C���g���ߝ� 2���V�h��ό�߰� ��Q���u�
���@� ��d��߈��)��M� ��������<�N��� r����%�����[��� �&��J��n� �3��i�� "�/X�|� �A�e�/�0/ �T/f/��//�/=/ �/�/s/?�/,?>?�/ b?�/�?�?'?�?K?�? �?�?O�?:O�?GOpO �?�O#O�O�OYO�O}O _$_�OH_�Ol_~__ �_1_�_U_�_�_�_ o �_DoVo�_zo	o�o�o ?o�oco�o
�o.�o R�o_��;� �q��*�<��`� �����%���I�ޏm� ����8�Ǐ\�n��� ��!���ȟW��{�� "���F�՟j���w��� /�įS��������� B�T��x������=��ҿa������,����$FILE_FR�SPRT  ��������A�MDONL�Y 1dU��� 
 �)MD�:_VDAEXTP.ZZZ3�俻����6%NO� Back fi�le ����eH��߫�@�	�M�v� ����)߾���_��߃� �*��N���r��� ��7���[������&� ��J�\��������� E���i�����4�� X��e��A� �w�0B�f����E�VISB�CKs�]���*.�VD��UFR�:\�ION\DOATA\�xU�Vision VD��/![/m/� �/{�/D/�/�/z/? �/3?E?�/i?�/�?? .?�?R?�?�?�?O�? AO�?ROwOO�O*O�O �O`O�O�O_�O�OO_ �Os_�_@_�_8_�_\_ �_o�_'o�_Ko]o�_��oo�o4oFo�o;�L�UI_CONFIoG eU��>�k $ �cx�{U�=Oas���y%p|x�o��� ��'��J�\�n��� ��)���ȏڏ���� ��4�F�X�j�|���%� ��ğ֟������0� B�T�f�x���!����� ү������,�>�P� b�t��������ο� �ϛ�(�:�L�^�p� ��Ϧϸ������υ� ��$�6�H�Z�l�ߐ� �ߴ������߁�� � 2�D�V�h��ߌ��� ������}�
��.�@� R�d������������ ��y�*<N` ��������u &8J�[� ����_��/ "/4/F/�j/|/�/�/ �/�/[/�/�/??0? B?�/f?x?�?�?�?�? W?�?�?OO,O>O�? bOtO�O�O�O�OSO�O �O__(_:_�O^_p_ �_�_�_=_�_�_�_ o o$o�_HoZolo~o�o �o9o�o�o�o�o  �oDVhz��5 ����
���@� R�d�v�����1���Џ�������Ro�bot Speed 10%�S�e�Pw���������x���  �$FLUI�_DATA f����ۑ�ɘRESUL�T 2gە�� �T�/w�izard/gu�ided/ste�ps/Expert��;�M�_�q����������˯ݯ�����Continue with G�ance��8�J�\� n���������ȿڿ��� ��-��ە�0 ����G�6ۑ��ps ψ� �ϬϾ��������� *�<�N����u߇ߙ� �߽���������)� ;�M海璪�M�/ϑ�:S�&c�rip&���ToolNum/NewFram&� �����#�5�G�Y�k��}������0x0 ��������'9�K]o���  A������S�c����imeUS/DST�;M_q���������Enabl��#/5/ G/Y/k/}/�/�/�/�/(�/�/�/����05?G?	24&�? �?�?�?�?�?�?	OOx-O?O�Dis/ uO�O�O�O�O�O�O�O@__)_;_M_5e��I?+?�_O?a?zon#P_�_�_oo+o�=oOoaoso�o�o��PST Paci�fic Stand��o�o�o�o" 4FXj|��� Ѳ��__�S��~ �Region� 3�E�W�i�{��������ÏՏ��Americav�!�3�E� W�i�{�������ß՟矦�qy?�1�C�����Editor ����������ϯ�����)�;�V� To�uch�`nel �p� (recommenn�)I����� ��Ŀֿ�����0�Bϭ|��#��ϗ�Y�>��acces��� �����"�4�F�X�j��|ߎ�M�Conn�ect to N?etwork���� ����
��.�@�R�d�v���x�i][P�y���^!���PIntroduct� 2�D�V�h�z������� ������Q���+ =Oas���� ���cRZU����1����/Safet �t������ �//(/:/��^/p/ �/�/�/�/�/�/�/ ? ?$?6?H?c?�? O�\�_�?�?�?OO /OAOSOeOwO�OH/�O �O�O�O�O__+_=_ O_a_s_�_�_V?h?z?��_�9#�?�6/current�_3oEo Woio{o�o�o�o�o�o��o��31-OCT�-18 01:42 PM�o$6H Zl~������W�T��_�_-��<9 �_gYeau��� ������ˏݏ����%�7�R�2018 A�j�|�������ğ֟������0�B� 
��������S�>gMonthD�ٯ ����!�3�E�W�i�8{�����10���� ο����(�:�L�@^�pςϔ�S���
q�d�ϙ>��gDaq *�<�N�`�r߄ߖߨ�0�����ߝ�31��� "�4�F�X�j�|���@��������Ϲ���p'�A���gHour� ���������������!3�g��bt ������� (:����{�>"O���inute@���//0/�B/T/f/x/�/��42 �/�/�/�/�/ ??$? 6?H?Z?l?~?�?O���*m�?=��gAM &O8OJO\OnO�O�O �O�O�O�O��O
__ ._@_R_d_v_�_�_�_P�_�_�_�r�r��p��?�?%o�&�6r�ippera�oo�lNum/Fraj�s��o�o�o�o�o �o�o�o#5LY k}������ ���1��?�?lv��8o)Ko]iActiveib<�ُ�����!�3�E�W�i�{�:
0xf������Ο�� ���(�:�L�^�p�����G�j���j�̯������Macro�e`s/New	�s ��-�?�Q�c�u�����𫿽�Ͽ��0x0 �	��-�?�Q�c�u� �ϙϫϽ����Ϡ�U����-ߟ,��	�Openno�ߓߥ� �����������#�� LY�k�}������ ��������1�H�Z���v���?�Summary8����� ����"4FXj |;�`����� �/ASew�C�M�ߩ����FRobotOp �/./@/R/d/v/�/ �/�/�/�/��/?? *?<?N?`?r?�?�?�? �?�?�?���#O���tutojo�g��Overview�?rO�O�O�O�O �O�O�O__&_�/J_ \_n_�_�_�_�_�_�_ �_�_o"o4o�?OOo�yo�"CO��electT1Modr� �o�o�o�o#5G Yk}<_���� ����1�C�U�g��y�8oJo\o��Џ�(��o��Enable�TeachPendant��$�6�H� Z�l�~�������Ɵ؟ ���� �2�D�V�h� z�������¯ԯ��Տȷ���$돩gJoinZ�gޯt����� ����ο����(� �L�^�pςϔϦϸ� ������ ��$������i�{��'?�UEr��_[���������� �/�A�S�e�w�6ϛ� �����������+� =�O�a�s���D�Vߠ�����ߢhHoldD�eadmanSwitch��1C Ugy����� ���	-?Qc u���������Ȳ�/ڍ ���aRe�setAlarm �l/~/�/�/�/�/�/ �/�/? ?�D?V?h? z?�?�?�?�?�?�?�? 
OO���IOsO�q!;/�a��_J1.O �O�O�O�O	__-_?_ Q_c_u_4?�_�_�_�_ �_�_oo)o;oMo_o qo0OBOTO�o�o:��OJ2-J6�o* <N`r���� ��_���&�8�J� \�n���������ȏ�o0�o�o���#�oQ�Car��g�y����� ����ӟ���	��� ?�Q�c�u��������� ϯ����)����D�n���&7���S��� Ϳ߿���'�9�K� ]�o�.��ϥϷ����� �����#�5�G�Y�k�@}�<�N���������I���_X~��!�3� E�W�i�{������ ��������/�A�S� e�w������������������O��_Y-Z��ew���� �����=O as������ �//������B/l/��o��_Rotation�߻/�/�/�/ ??'?9?K?]?o?. �?�?�?�?�?�?�?O #O5OGOYOkO*/</N/0p/�O���/onQ_ !_3_E_W_i_{_�_�_ �_�_�?�_�_oo/o AoSoeowo�o�o�o�o��k�O�O�o- ��OI�LastScreen�o`r� �������� �_8�J�\�n������� ��ȏڏ����{O�o��o=�g�--/ugr�ipper��Ma�croNum��CloseUse"� ��ӟ���	��-�?�Q�c�"�2q����� ��ͯ߯���'�9�K�]�o�-�
*�m��a�M����߃���Set?Methodt�� �+�=�O�a�sυϗ���ϻ�&�Dire�ct entry� of EOAT data���� '�9�K�]�o߁ߓߥ�$����-���������w/ٿ�trai�ghtOffset��`�r�����@��������+�A� Tool�K�]� o��������������� ����9�����X�M%+I��/�� ��� 2DV|h+�50.0� m������/@/)/;/M/_/p-��iBH  M�/q��Yp/	??-??? Q?c?u?�?�?�?�?|85��?�?OO0O BOTOfOxO�O�O�O�O/�*��/_�/�/�Z�O]_o_�_�_�_�_@�_�_�_�_o,��? :oLo^opo�o�o�o�o �o�o�o �O[-���OWZ)'_��Ro�tation�wW ������!�p3�E�W�o18� ������Ə؏����� �2�D�V�h�'eyC�4G��k}�onPl�	��-�?�Q�c�`u�������j�-�? �����+�=�O�a��s���������z�<
����������ӟ�R��]�oρϓϥϷ� �������Ͼ�(o5�G� Y�k�}ߏߡ߳����� �����̿6��R�[�"#�5�tp3Zdir/Tp3z� �����������(� :�L�^�߂������� ������ $6H�Z�+�=�c�#P+�w�5�Measur�ement/StraighJ_ );M_q��� f�x���//%/7/ I/[/m//�/�/�/t����/��/We��Nums/New53s�/[?m??�?��?�?�?�?�?�?l�0x�4OFOXOjO|O �O�O�O�O�O�O�O_�s��/-Y�/O_i�.�?1<Tool53Use_�_�_�_�_�_�oo0oBoToo�1 ao�o�o�o�o�o�o�o�);M_s�
#_�$=_�a_s_1<Part�_��!� 3�E�W�i�{�������pb2��ۏ����#� 5�G�Y�k�}�������Dr�)��e�(�17s/G� 53��T� f�x���������ү�<����12�0� B�T�f�x����������ҿ�����/�A@��/I�g�)�-�Pa�yload1Cm B��Ϻ����������&�8�J�\��EO�AT w/o p �p]ߏߡ߳������߀����1�C�U�� �5_{���y��y`� ��� �2�D�V�h�z� �������������
 .@Rdv�� ���/;��_����2��N`r���@����/��q�ithy�3/E/W/i/ {/�/�/�/�/�/�/�/@d����&?P?��&�)Advanced?�?�?�?�?�?�?�O O2ODOVO��0x���O�O�O�O�O�O �O�O_"_4_F_X_��A?-?w_�_��%k?�)Mass/Center�Q\_�_o o+o=oOoaoso�o�o �o���o�o�o' 9K]o�����v_���_�_ss ��M�_�q������� ��ˏݏo�o%�7� I�[�m��������ǟ ٟ������B��),�)Gt0c�R-�X�����ȯگ��� �"�4�F���|��� ����Ŀֿ����� 0�B�T��%�7���[�m��sYX���
�� .�@�R�d�v߈ߚ�Y� k���������*�<� N�`�r����g�y�`���������sZ�� L�^�p����������� �����߿�$6HZ l~������@�������A�.� !�#!-������� ��//1/C/ y/�/�/�/�/�/�/�/ 	??-???Q?"40�?Xj|rt���? OO+O=OOOaOsO�O �OV/h/�O�O�O__ '_9_K_]_o_�_�_�_�d?v?�?�_�?�?�?rt:�Io[omoo�o�o �o�o�o�o�O�O!3 EWi{���� ����_�_�_>���lTCPVeri�fy/x�Method�������ҏ������,�>��lD�irect EntryM�~������� Ɵ؟���� �2�D�� x�m�-����Z'_�q�fy�����  �2�D�V�h�z�����	p50ȿڿ� ���"�4�F�X�j�|�0�Ϡ����BH+��� ����ǯ�?>�P�b�t� �ߘߪ߼������߱�85���.�@�R�d� v��������������ʪ��5���	�� 8o�������������� "4F	j|� ������ 0B�/�)��I�[�m�fyWL��/ ///A/S/e/w/�/�/ �18���/�/ �/�/??0?B?T?f?`x?�?�?[�C4{�?���P�?;OMO _OqO�O�O�O�O�O�O�O��-
�_)_;_M_ __q_�_�_�_�_�_�_x�_�?l�����?3o�?Ou�R�_�o�o �o�o�o�o�o1 CZgy���� ���	��-�?��_�hz��Fm*WoiofyMeanH���� 
��.�@�R�d�v����/*����Ɵ؟��� � �2�D�V�h�z���@K�]���y�ۯIj)����πax��9�K�]� o���������ɿۿ�� ���#�5�G�Y�k�}� �ϡϳ������Ϩ���̯.�Hk"���In�troductioԏ�ߗߩ߻����� ����'�9�Put�X� j�|����������@����0�B�Op���a���Qb S�fi�le/backu�p�device F������� 2D�Vhz�OvFr�ont Pane�l USB (UD1)���� );M_q��_   Op�Op!��s��Gl%�����irectories�1/C/U/g/y/��/�/�/�/�/�/Tq�� :\\BKUP�_28-NOV-�18_12-04-58\\�/-??? Q?c?u?�?�?�?�?�?��?�\���6O��q!���WAdef�? �O�O�O�O�O�O�O�Op_#_5_PuSy�m B�� ZRc_u_ �_�_�_�_�_�_�_o0o)o;o���O�yo�o�$OO��Summary/S] �o�o�o1CU gy������ �	��-�?�Q�c�u������Ojo�oޏ���S�crea�r;og�Groa_$� 6�H�Z�l�~�������xƟ؟�0x2� ��1�C�U�g�y����������ӯ�  �O��Ï%��o�o�l1 诀�������ȿڿ� ���"�4��/	??|� �Ϡϲ���������� �0�B߭��u߇�I�[�S��������	�� -�?�Q�c�u��J_� ����������)�;� M�_�q�����T�f߈� ��LO�ߛ�%7I[ m������ ���,>Pb t��������  O�� /*/��"��aE�ress�z/�/ �/�/�/�/�/�/
?? .?�R?d?v?�?�?�? �?�?�?�?OO*O:LA�/UOO��,G/Y-`&6:O�O�O�O_� _2_D_V_h_z_�107�_�_�_�_�_�_ oo/oAoSoeowo�o  ��]O�o�o�O �O�L�_+=Oas�������94���(�:�L�^� p���������ʏ܏�o��o�o!��o�os8 ����������ȟڟ�����"��|	SYS�UIF.SV��AME.TP1�h�z� ������¯ԯ���
� �.��/��s���H? ����˿ݿ���%� 7�I�[�m��B?�ϵ� ���������!�3�E� W�i�{ߢ��у�]��� �ߓ���
��.�@�R� d�v�������� ����*�<�N�`�r� �������������߯� ��#��J\n�� ������" ��FXj|��� ����//���� u/7�/�/�/�/ �/�/??,?>?P?b? t?3�?�?�?�?�?�? OO(O:OLO^OpO�O�A/S/e/�O�&C�g�uidedV�NetDone�O_&_ 8_J_\_n_�_�_�_�_ �_�?�_�_o"o4oFo Xojo|o�o�o�o�o�o�I�I��O�o=��C�networkV�Port�ofx ����������5�Qq 1 (?CD38A))�\� n���������ȏڏ�p���"�H� �`��`%i��O=�s/method ,���Ο�����(��:�L�^�p��ZManual}�����̯ ޯ���&�8�J�\�n�-�?���ay�[����,��MqSummary���#�5�G� Y�k�}Ϗϡϳ����_ ������1�C�U�g� yߋߝ߯�����F��o������ݿGw�@TesTd�v����� ����������<�N� `�r������������� ��&����	�k�& 7�Mqsett?ingsp1*� ���(:L ^p/������ � //$/6/H/Z/l/@+=O�/�/�B�>MqIntro~/? ?/?A?S?e?w?�?�? �?�?~�?�?OO+O =OOOaOsO�O�O�O�O@�O�o�/�/_�%�/>�/name�Oi_ {_�_�_�_�_�_�_�_�oo�1ROBOT!oKo]ooo�o�o�o��o�o�o�o�o# �G_�Oa{&3_E\ipad����� ���)�;�M�_�q���1192.16?8.1.40u��� ��ʏ܏� ��$�6� H�Z�l�+=O��ßs�'�E\sub?� x��%�7�I�[�m��𑯣���ǯ �255.ݥ������ 0�B�T�f�x������� ���������ٟC^?router̿g� yϋϝϯ��������� 	���??�Q�c�u߇� �߽߫��������� ֿ���\�z$/�E\mac ��������  ��$�6�H�Z�l�+��00:e��4:�41:8b:b9 q����������� %7I[m,�n�P� ��+0���/ ASew���� *���//+/=/O/�a/s/�/�/�/�/�H � ���/?�6?H? Z?l?~?�?�?�?�?�? �?�?O�2ODOVOhO zO�O�O�O�O�O�O�O 
_�/�/�/�/a_#?�_ �_�_�_�_�_�_oo *o<oNo`oO�o�o�o �o�o�o�o&8 J\n-_?_Q_�u_ ����"�4�F�X� j�|�������qo֏� ����0�B�T�f�x� �������������x#���NetT�est/ipaddß[�m���������ǯٯ����΃1�92.168.1.40�F�X�j�|� ������Ŀֿ����`{��Q�c��&'��9�linkstatϲ������������0�B�T�f�р	ConnecteI� �ߨߺ��������� &�8�J�\��-�?ω���!�!{ύ�url l���%�7�I�[�m���������̅http://)����� 1CUgy� ��n����� -?Qcu��� ����/ȏ)/;/ M/_/q/�/�/�/�/�/@�/�/?ğ֟�� W?~?�?�?�?�?�? �?�?O O2ODOVO/ zO�O�O�O�O�O�O�O 
__._@_R_d_#?5? G?�_k?�_�_�_oo *o<oNo`oro�o�o�o gO�o�o�o&8 J\n����u_ ��_��_"�4�F�X� j�|�������ď֏� ����0�B�T�f�x� ��������ҟ���� �)��M��t����� ����ί����(� :�L�^���������� ʿܿ� ��$�6�H� Z��{�=���a�c��� ����� �2�D�V�h� zߌߞ߰�o������� 
��.�@�R�d�v�� ���k��������� *�<�N�`�r������� ����������&8 J\n����� ��������+U �|������ �//0/B/T/x/ �/�/�/�/�/�/�/? ?,?>?P?Y3}? �?i�?�?�?OO(O :OLO^OpO�O�O�Oe/ �O�O�O __$_6_H_ Z_l_~_�_�_a?s?�? �?�_�? o2oDoVoho zo�o�o�o�o�o�o�o �O.@Rdv� ��������_ �_�_K�or������� ��̏ޏ����&�8� J�	n���������ȟ ڟ����"�4�F�X� �)�;���_�į֯� ����0�B�T�f�x� ����[���ҿ���� �,�>�P�b�tφϘ� ��i��ύ��ϱ��(� :�L�^�p߂ߔߦ߸� ������ ��$�6�H� Z�l�~�������� ��������A��h� z��������������� 
.@R�v� ������ *<N�o1��U� W���//&/8/ J/\/n/�/�/�/c�/ �/�/�/?"?4?F?X? j?|?�?�?_�?��?��?�$FMR2_�GRP 1h�5�� ��C4  B�0	� �07OIL4@E�� F@ _Bǂ5UkE�*4@J���NJk�I'�PKHu��IP��sF!��wM?ǀ  �O�<4@9��<9�8�96C'6<�,5��wMAg�  �O[BH1C�B�-@,PQ@�3]37R�33�<3DxY_j]4@@UUUZ�@5P�PwM�)>u.��>*��<����wM=[�B=����=|	<��K�<�q�=��m�N��8��x	7H<8��^6�Hc7��x�_ ok_oVoAo�zoeo�o�'B_CF�G iKT ��o�o�o�kNO� J209693   �m�RM_CHKTYP  
A�0"@$@��0AROM_p_MsINep�3���pu�PPX@SSB�c�j�5 5F��5�s���e�TP_DEF_O/W  �4"C��IRCOMdp���$GENOVRD�_DO�v�!C�T[HR�v d`�dI�o_ENB5� I��RAVCCk�w�p �WEG|� Ga� G(�� I�W�I�x�JM+ȃo���}F�$�GZ �V��OU@qLKqqGH�GE<�p��O��E�����㟵3C�  D����-�R=�A�W*�B�)�pJI�����SMTC�r��&@�p��$H�APTIC_CNoT 2s�5��}
�r��@���2A,@���%�7��I�[�����FEAT�  ͦ��� <�s���uq����ɻ��O3STŠ�`1tI�p���/ 	��&�����&+ϯ)eG�xϊϜϮϮ* f�������8�9����	anonymous<�j�|ߎߠ߲� ������2�T��� C�U�g�y��ϝ���� �����>�P�-�?�Q� c�u������������� (�);M��q �������$� %7I������� �������/V  /E/W/i/{/��/� �/�/�/�/?Rdv ��/d?��?�?�?�? �?*/OO+O=OOOr? �/�/�O�O�O�O�O&? 8?J?�O^OK_�?o_�_ �_�_�_b_�_�_�_o 4_5o|OYoko}o�o�o �O�O__�o2oT_1 CUgy�_��� ��>oPo-�?�Q� c�u��o�o�o�o�� (��)�;�M��q� ������ʏ�������%�7�n�ݱEȠ1�u��  P!\˟��  Z�w� ����د������ �� ,��U�z�=���a�¿ ��濩�
�Ϳ߿@�� d�'ψ�KϬ�oρ��� �����*���N��G� ��sߨ�k��ߏ��߳� ����%�J��n�1�� U��y���������4���X��QUI�CC0e�A�!1�92.168.1.41��s�����R��v�2����T!ROUTERU�1C�!PCJsOG��!���0.10~�s�CA�MPRT����1�RTn 2��Y�NAME !~f�!ROBO��S_CFG 1�tf� ��Auto-st�arted��FTP��,!����W/ �{/�/�/�/�/`��/ �/??@/.?�/e?w? �?�?�?~�//)/O =?_/ONO`OrO�OK? �O�O�O�O�OO�O&_ 8_J_\_n_�_������ ���O�_3Oo"o4oFo Xo_|o�o�o�o�o�_ io�o0BT�_ �_�_��o�o�� ���o>�P�b�t��� �+���Ώ����� ]o��������� ��ʟܟ��$�6� H�Z�}���������Ư د�1�C�U�2�i�V� ��z�������w�m�� ��
��?�@�ӿd�v� �ϚϬ����)�+� ��_�<�N�`�r߄�K� �ߺ�������ߕ�&� 8�J�\�n�������� ������3��"�4�F� X��|����������� i���0B��_ERR v��RbPDUSIZW  ��^��y�>�WRD ?�����  guest������,�S�CDMNGRP �2w�| C������4��Kq� 	P01.0�1 8�� ������  �    
=�� ������*���u�������ù�/X�&/'2����U��ఱe�����������O�m P���y1/ؑ/�!��d���|�J_GROU\Uxq	s>	T��69QUPD � ��y	4E0T�Y�0qd TT�P_AUTH 1�yq <!i?Pendan8�>�A�=�2!K?AREL:*�?�?�=KC�?�? O�0�VISION SET0^O5O�7�� cO�O!�O�O�O�O_��O�OD__-_}4C?TRL zq���X
�0^FF�F9E3R_��F�RS:DEFAU�LT�\FAN�UC Web Server���Pb �1��uL.ne\>oV_�ro�o\WR_CONFIG {`� o�_bIDL_CPU_PC�P���B����` ?w���cMIN�l��`�{PIGNR_IOk���w�`�NPT_SIM_�DO0v:{STA�L_SCRN0v ��S8INTPMODNTOLrw:{aRTYQx�a?vR@�0�ENBrwR2�dO�LNK 1|q � ��&�8�J�\�n�>�rMASTE/pJ?��qSLAVE �}q�tSRAMC�ACHE�����1O�_CFGΏ��UO�h0��r_CMT_�OP�P2ru
$�YC�L͏!��P_ASG� 1~`�
  p�������ɟ۟��� �#�5�G�Y�k�}�x��f�NUM�u	
��IPˏ݇RTRY_CN/�!�nqb1���y ��낃��� <�� �`R�CA_ACC 2��;  M|`��T�� ��� 27� 6�Q����p��� ��r� ����bU�oBUF0�2�;�= ]@u1
�8j�]`u4�3]]�u1��m�]�u2�q`�]�u1��gi]�u3��`�^ u1��hp^ u1 �"�^�-�`+�� �@T�^�+��u�2Z1^�u�1�qY_ u�3�^i_*��j!_@c�"_�_:��l�`� t��b`� u2�h�`�@u2�_�`�:�
9j�`�u�3be�`�u�4{b�`�u�2�eA`�?�pXXZ�-��Y"���*�Y��-�2EY:�Y���J�Y�T����Z��Z*�Z2�}Z:��X�Z�_xq�ZJ�Z��UZ��[��[*�[2��[:�[��[�u3� U![���s�[�u4"k�R�\��\��y�Y�\�]�\`u�7?U�\����t�\r��[i�\�u4,m}\Z� Z1]"���m�]��`й2ݿ�+���u4 ����
�������u�P!�+�)�.� ��9�.��I�.�R��� Y�+�a�&�i�f�r�n�C��tӈ������� ����&���������`��+�����3� �������������� �+�	��3���C� )��S�9��c�I�N� 3�Y�N�C�i�N�r�&� y�N����+������і��u7���� &�ю�c����ғ�й3��ﳰ!����� �� �!!�/*�8� /:�H�/J�X�/�� h�o<q�oL��� ���� ������ �������!����� <������� �� l	��!� 1�@�lI�X�W a�p�Wr�W$�Ѱ! �Ә��ї�� ��Зl���R��2�=�Q)�%� <� %$(!2r�R�HISڲ�;� �p� 2018-11-28�&� �( 2r( *{$ {$({$0{$m"z( @�Q; H�1�9 � X�"!5 `uQ8 �`�  7 �	���/??(=M{�`b(�r/�/�/�*�&"� &"]B( � �!T� &"hW4pW4xW4��W3��( �W4��W4��$��$�W4��W4��1( Mz<:6�J?\?n?�.�"�  + ��"�8�"�?�3�4 �8�2�8�2�4Q�0�2Ny<:5&O 8OJO�?�?�2&"�?�C �0�"�0�"���2�?%#�0&"�?Dx<:_�_*_<_N_  : f_�"�0=b�O�_�_�_Mw<:.�_�_oo*l� �"� "�!�@�"vT�<io{o�oIv<:��o�o �o�o*o`_�O<N`�r;+��L/^/�z(!d ����p���p���p����p��m ��� ��� 0������� ��� � ��(?�*�<�*?<?�� ����͏� ~��}�� ~�
�~��0~��P~����~�*�~��0~��0(!c �0~�J�~�@~�@~� Oq���������� !r
� 9�0`۟����d�-��ON�`�r��� ��̟��̯ޯ��8� �_*�<�N�`�r����������P˿ݿ7��o ��*�<�N�`�rτ� ���Ϻ�8������� �*�<�N�`�r߄ߖ����=)��q����y�Z�	!���� ��(���0��8��@ ���	!H ��	!P� �z	!X �j�	!` �u� �q)6�H�Z�l�Z�l�S������� ��U(��0��8��@���H��P��X �At���h��p ��x	� ��	!����� �U�	!�������c�`��;��y����~} }(}0z}8}@ � �ۏ����q��'���p�x� �Y����� ���� �M<�oD���#�`����y}�1��ZY Y(Y0�Y8Y@YHYP�YX }��h� }�TM���~�}U�}�}�}�}��}�`~�yx����6#5$ 5$(�5$05$85$@5$H�5$P x��z��#h zE|M}I�#��$U��$�Y�Y�Y5�Y�Y�`Z�Ϧ�yl��34 �4(40484@:4H4P l*�p[p�sg��v��T 6#x5$�5$�5$U�5$�5$�5$�5$5�5$�5$�`6#��@??*?<?N:�2X�4U`�4h�4p�4x�4U��4��4��4��4U��4��4��4��4�`�3b�I_CF�G 2��� H�
Cycle �Time�qB�usyy�Idyl�B�Dminv�>+�Up�F�A�Read�G�Dow X�O\`Q��CCount�A	Num �B�C!y��|]�p�!b�SDT�_ISOLC  ����(p�Aw��$�J23_DSP_?ENB  �[�BJINC ��]ԗs�PA��?�=�?��<#�
�Qi:�o &a?oQo�q<oyo�WOBPR�OC�S�r(�f�aG�_GROUP 1퇳[��<� � aw��o�o?"y��_�pQ4Y k}<����y��io�iG_IN_�AUTO�dj�PP�OSRE�o�fKA�NJI_MASK�=�%�KARELMON ���_+ry���Ǐُ��� ��s��B�����S+t�:��TKCwL_L�NUM�P�T�$KEYLOGOGINGQ����/���U�PLANGUA_GE ������DEFAUgLT ɑ�QLD�A�-��TYX�Uϑ�GԒ�ڙWR �+q7�o���� ��+p'��y��+p;�+p�� ;���
r�(UT1:\��� ������ ůܯ����$�1�C��l�(�����VLN_DISP ��_�	X31�OCTO	L�߱D�Ra���GBOOK ���dc�Qf�f�3� ��W�i�{ύϟϱ�`��!�S�ɯ�	�@��a���,�Q��_BUFF 2���[ -ߺ� b�2��~�W�߬��� �������E�<�N� {�r�������������CF�DCS �ڝb���y��Es��������"�IO 2�ڛ �@���@�P�����*: L^r����� ��$6JZ�l~���ER_ITM�^d���/ !/3/E/W/i/{/�/�/ �/�/�/�/�/??/?pA?S?���SEVQ���]�TYP�^���?�?�?b=6�RS�Tr� �SCRN__FL 2����P�S�SOeOwO�O�O�O��O�?TP���_�2>�NGNAM�TL�ܻ��UPS��GI�@?��U.Q_L�OAD�`G %��J%	SCAN_�SLO@w_�XMA?XUALRMo�?������U
�R4Q_PR9T?� �a�PC�����υ݆]��P�`P 2��[k �r�	�Af`+2���_ߴFbro]o oo�o���o�o�o�o�o �o1U@y�n �����	��-� �Q�c�F���r����� ���̏���)�;�� _�J���f�x�����ݟ ȟ����7�"�[�>� P���|�����ٯ�ί ���3��(�i�T��� x���ÿ���ҿ��  �A�,�e�Pωϛ�~��Ϫ��όWDBGDEF ��E�Q�Q�����_LDXDI�SAP�K��MEM�O_APPE ?=�K
 ��� l�~ߐߢߴ�������~�PISC 1��I�P���7�Ad�M���φ�q����_M?STR �{=��SCD 1�[ݠ �����@�+�d�O��� s������������� *:`K�o� ������& J5nY�}�� ���/�4//X/ C/U/�/y/�/�/�/�/ �/�/
?0??T???x? c?�?�?�?�?�?�?�? OO>O)ObOMOrO�O �O�O�O�O�O_�O(_���MKCFG ����_�SLTAR�M_OR�,geR�9`&RФ_�T�PMEgTPU7лc�����ND#`ADCOLx�U��^CMNT�_ �UFN`o�WFSTLI(og�� ���{n�S�Q�o|�d�UPOSCFIg=nPRPMo�i�ST�P1��� {4@P<#�
q #Qu'5w57I �m����� �-��!�c�E�W�������QSING_C�HK  +o$M/ODAQ�S��c[�eYωDEV }	��	MC:sW>ւHSIZE7�P��ӅTASK �%��%$1234?56789 t����чTRIG 1�.�� l��%��џ�S����ޟ��V�YP�A���҃EM_?INF 1��W��`)AT&�FV0E0��)�g�E0V1&A�3&B1&D2&�S0&C1S0=>n�)ATZ�ӯ��Hׯ�����'���A/�W��{�b����� e�ֿ��������0� �Tϋ�xϊ�=���i� ������߻�Ϳ>�� �φߑ�Kϼ����� �ߥ����:�!�^�p� #ߔ�G�Y�k�}���� �I�#�H���l�'��� ������y�������� ��DV	�z���Y c�����.�� R);�_� �/�*/�;/`/�G/�/l^ONITO�Rd`G ?�  � 	EXEC�1S�"2�(3�(4��(5�(���&7�(8
�(9S�"N24�" 24�"24�"24�"24�" 24224224 224,2�232982E82Q82�]82i82u82�82��82�82�83983�E83�"ӁR_GRP_SV 1�T�� (��������?l��fy���ү��6LϿ�$�-^�_D�#"D��CION_D�BQP��Q�@�̗P�@bT�D��@�G��@P̛ez N � '`	O��L��@�bU-u�d1-�C_U_g_�QP�L_NAME �!ke�P�!M�-10iA/12�, HandlingTool �S�wTRR2KA 1�� l<�QP
l d�b�_ �_oo%o7oIo[omo o�o�o�o�o�o�o�o@!3EW��2�_ ������� ��$���<qN�`�r� ��������̏ޏ�����oX2RrR=�N�
=�r�rTPa����� ԟ���
��.�@�R� d�v�������{���� ����*�<�N�`�r� ��������̿޿𿿯 ѯ&�8�J�\�nπϒ� �϶����������"��4�F� G| Gz  G��@<rUg@  �s߅�rRdo�WФ߶ݚ��� ��X�K�mZ���.��Q�T� A�l�b� t��������g@� h��rRA�	`V��P�b�t�3�:�o�A�R�������� A�  ��;� @7�U&0�R�S��Y�P>�, �� z"�Pe  @D7�  x?�~d�?rP�rQA/��xx+�oX;�	l��	 �x7J� �b@
P��  �< ��� � ��g@K��K ��K�=*�J���J���J9���E��Gg@@�t��@{S�`�(�El�#2�=�N����I��T;g�a����.Q+�*  �´  �� �>ʾ��~rQ?z����rQ�g�Jm�� /�"�##��.	�5��  {  �@X ��@�  ���@�p&���/1	�'� � �"�I� �  y���/:�È�/?È=����%4j�	��_ �n3��H/j"?m[j�6./Qz?  '��6]�@2��_@���@�@��@�C�CPC��@ C�C�C<��A�Ac �W  �B@�0
.BP(A�����1PErQD`���uO�7�O�O�O�O�@��( �� -��"�E�1�EnqrQ����  rP�р?�ff��._@_�OC -�u_�[58=0��_�Z>�!��,(=0�UP�X�I���^B3?��=0x=0���<
6b<�߈;܍�<��ê<���<�^�MoW��2:8��
j���?fff�?c ?&�`�@��.�b�J<?�;\��bN\�:9�2 �a�,��o~�ong �__4XC|g ������:8�eF���6��Z��o`{��iM���I�F�a��F�=2GI FU҃D��������PO�:�s�HL=3B>�A{�_����󛵟 �q�7���^�џ����8����N��b��M_A @|t��p��1��.�g���A���9O=5CT���P�������'���:9Đ���:�Cz u�CH7�$�Ĕy� ���@I܀��(hA� �A�LffA>�v??�$�?��Q+�°u�æ�)��	ff��t��#�E��g\)�=1@�33C|������<������G�B����L�B2�.����	b�+H�ۛG���!G��WHƥ�CE���C�+��<�I۩I��5�HgJF��y�E��RC��j=|�
�pI����G��`H����E<YD0;����������6� !�Z�E�~�i�{��� �������� ��D�V� A�z�e����������� ����@+dO �s����� �*N9K�o ������/&/ /J/5/n/Y/�/}/�/ �/�/�/�/?�/4?? X?C?|?�?y?�?�?�? �?�?�?O	OOTO���(�����ob�y��E@E��xO<�O��3�8��O�O��4Mgs�O�O��ϴVwQ�O_4p?�+4�](](Y�h_V_�_z_�_�\ٵPHbP�^����o^O`oAo,oeoPkRko�ro�o�o�o�o�o  )P��o�o/S>�wo����{����$�J�8� �R�AS�e������������  2 G���Gz��G�膞�B�������t�C喚�@����8�����<Z8��p8�u8�T�@�T��6��J�����sEQ�sI���ܶ�a��(������,���?��W�@@��؄�����oq��ܾ
 :�������ӯ� ��	��-�?�Q�c�u������w� ���KX��ʘ�$MR_�COM ��X���n�P4�T�&%% 23�45678901���� ���#���#�E�#�#�
�Ǔ�not ?sent *o�#��?�W�UTE�STFECSALMG�`egʚE�d��`k�C������P��P#���=��������� 9UD1:\�maintena�nces.xml��\�  z���DEFAULT�Ŝ��GRP 2�|˺�p�  �l���#�  �%�1st mec�hanical �check�#������ �	�l� �P̚4�F�X�j�{������controller�Ԫ�����m�%�����0���cM��j�#�"8��!#����l�������������@�%C ��0�T�����������C��g�e��. batt�ery�Dl�	 qFXj|��	���dui��able^�  Dp�֒��5
//./@/�R/���greaYs�@�f��#-#��!�/l���/�/�/h??��
�oiJ��/�/�/�/�?�?�?�?�?���
�#���C<#�"A)Ol�
�?VOhOzO�O�O�!t�O!O�EO_�,_>_P_b_��Ov�erhauc��L��R x#��Q�_l�	_�_�_oo&o#�$�_No��ͳ˸vo v �_�o�o�o�o�o:o ^opo�oCi{�� � �$6H�/� A�S�e��v������ ������+�z�O� a�����ԏ����͟ߟ �@��d�v�K���o� ���������ۯ*�<� �`�5�G�Y�k�}�̯ ����׿&����� 1�Cϒ�g϶�ȿ��� ��������	�X�-�|� �Ϡϲχߙ߽߫��� ���B�T�f�'�M�_� q����߹���,� ��%�7�I���Z�� ������������� ^�3E��i���� ���$�HZ/ ~Sew����  �D/+/=/O/ a/��/���/
/�/ �/??'?v/K?�/�/ �?�/�?�?�?�?�?<? O`?r?�?�?kO}O�O �O�OO�O&O8OJO_ 1_C_U_g_y_�O�_�O �O_�_�_	oo-o?o�T	 @@omoo�_ �o�_�i�o�o�o�o * `6Hr� ~�����&����\�n�D�N� ���Q?� Zc  �o��ӏ參V���$��6��X*V�** ~�|��p��������p�ҟ������ �_�Sm��Y�k�}�?� ����ů�!�3���� 1�C���O�y������ ��_����	�S�ݿ?� Q�cϭ���ѿoϽ��� �ϣ���)�sυσU��$MR_HI_ST 2�|����� 
 \�R$ �23456789C01�ߘ�Y�P���9�_������_I� [�m�$�6�����~� �����!���E���i� {�2���V��������� ��/��S
w� @�d�����l�SKCFMAPw  |���U�� � �ONREL  �d�8i�SKEXCFENBjq
6�FNC��|JOGOVLI�Mjd���!KE�Yj��_P�ANi��!RU�N��SFSP�DTYP�u S�IGNj|T1M�OT�y!_C�E_GRP 1�|�8��X`��/ ��/�/e��/)?�/M? _??�?:?�?�?p?�? �?�?O�?7OIO0OmO $O�O�O�O�O~O�O�O �O!_�O_W__{_^��D _THRSHD�  �F@ ��QZ_EDIT�g$2�STCOM_�CFG 1�.���_oo 
�Q_/ARC_�dյ�T_MN_MOD�Eg&�UAP�_CPLDo�NO�CHECK ?^.  �o �o�o�o%7I [m����S�NO_WAIT_�Lf'�W� ODRD�SPCci&�OFFSET_CAR�P��o9�DISF�7�S;_A^`ARKg'�Y�OPEN_FIL�Ee�i!"a�V:`OPTION_IO�����M_PRG %.%$Y�����WO����'�FB��9�=T�� ; E�S���S�	 ��S���s���RG_DSBL'  x�8>T���VORIENTT�Oi�RC�H7A� 7�UT_SIM�_DŇ5���V~�LCT �.��TL�"a>����_�PEXf`h�W�RA-Tfg d�W�>��UP �"����M����˯������$PARAM2�#�� }l�
l dr_ D�V�h�z�������¿ Կ���
��.�@�R�@d�vψϚϬϽ23� ���� ��$�6�H�Z�l�~��<�Ϩߺ��� ������&�8�J�\� n�4^�<��	栨����P����
��.� @�R�d�v��������� ����������<N `r������ �&8J+ �������� /"/4/F/X/j/|/�/2�.olW��/�-Q�pT�/>�/2?@7��-�-q_�?n?�?Z7 ���7�?�?�?�?�?O�"ODO�0,�gOwL�r�5	`�?�O�O�O�A:�o��O�O_|"_�0A�  9Y �?Z_�<G�|_�X���O��1� ˌ� ��(��B�, ���р�P �@D�  �Q?���S�Q?�p�Q�qD��R�Q���x;�	�l�R	 ��xJ0`��F�G�'` �<w �F`� �Lb�NPH(��H3k�7HSM5G�2�2G���GNɁ3i\���/�o�lNPC%f�a搿a��c�Q��oKS�����4
�`>�`�`u��o�o��<B_����=j�q�tq. flr�Q�sNW�Y�oNR�b�{  �@ᐊƀ�  �7���vN_�JU	'� � 
��I� �  ��FUHV=���P.�@��s�Q	:P��p�nb�⾦����D�뎒u_�~HXN�؏  '����a�}C�C�@ C#p�C'pC+����� � �A�pzhB�`��xjv�J��pB�򐆑9_+[S����Rz G_џ0�����+����( �� -�O�K�[���&����Y����!�?�ffQ?�����0� �@ӯ��8����	�>O�l�Q�	(��7�P@�[�=a6c�6d��?����x�����<
6b<�߈;܍�<��ê<���<�^�no����R�����R
���R6P?ff�f?�p?&��@��.���J<?w�\��N\��� R���m��U>��W]� ̷"d����}϶ϡ��� ������"�4��X�j� Aߎ�y߲�)�K�Mϫ����F�  GF����GI FU 0��S�>�w�b�t��H����|�L[��@A�� ���l_?�Q��	o�� ���߼�/�����α��b����A @|��k���z0����AA�����YEC��t�&?��EL�pym��D�ȘC�PF�CH���_�_�^!@I���(�hA� �AL�ffA>�v?��$�?�C�	z���u�æ�)��	ff��t��s#�{�=+g\)YA�@�33C|������<��:.G�B����L�B2�.?����	t�	z�H�ۛG��!�G��WHƥC�E���C�+��}I۩I�5��HgJF�y��E��RC�j�=�.
�pI����G��`H��E<YD0 �:?L?7?p?[?�?? �?�?�?�?�?O�?6O !OZOEO~OiO�O�O�O �O�O�O�O __D_/_ A_z_e_�_�_�_�_�_ �_
ooo@o+odoOo �oso�o�o�o�o�o �o*N9r�o �������� �J�5�n�Y���}��� ��ڏ�׏���4���X�C�|�g�y�����(Ξ���[�m���<敞���֟�>!3�8���>!�4Mgs.�@�>!��VwQZ�l�4p�+4�]����Ư@���د���7P��	P@�_�\�i���u�0����ÿ��Rɿп`	����?�*�  ���B�Tύ�xϱϜ����|�N����,�� 2�<�r�`߂ߨߖ�< ������������A��O�  2 GvYGz;'G��>&�B�� �� �C���@�������������=��I�[�m�����>#?���@U@a*��> > �9�> :
  ����1CUg y������<*��� ��*�X�����$PARAM�_MENU ?���� � DEFP�ULSEa+	W�AITTMOUT�IRCV\ �SHELL_W�RK.$CUR_oSTYLG��OPT��PTB���C�R_DECSNT1����/ "/K/F/X/j/�/�/�/��/�/�/�/�/#?S�SREL_ID � ��Z��25US�E_PROG �%-%?�?33CC�R`D2Z�5�7_H�OST !-!�4�?�:TQ��?�3ļ?�1�31O�;_TGIME^D6�5?GDEBUGB0-�33GINP_FL'MSKZO�IT尚O��EPGA�@ yL�8��KCH�O�HTY+PE*6�?? N_w_r_�_�_�_�_�_ �_ooo&oOoJo\o no�o�o�o�o�o�o�o �o'"4Foj|��������EW�ORD ?	-
? 	PRv@ֳ�MAI�ײSU�:�TE@ֳ�xs	�G�COLԵ�c����FTRACE�CTL 1����7 ��� }�Y� � ����\�Y�ۄ��DT �Q��� �ŀD� � WȁU�	�
��U����TD0������7�8�0��Ё�؁����@�@�������� �"�4�F�X�j�|��� ����ğ֟����� 0�B�T�f�x������� ��ү�����,�>� P�b�t���������ο ����(�:�L�^� pςϔϦϸ�������  ��$�6�H�Z�l�~� �ߢߴ����������  �2�D�V�h������	�\w�\:V����\��\��\'�\�/�\7�\��\��\���\��\��\��\���\��\��\�\*�\_�\g�\o�R� d�v������������� ��*<N`r ������� &8J\n�� ������/"/ 4/F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?f?x?�?�?�?�?�? �?�?OO,O>OPObO tE�O�O�O�O�OJ�qE �_�_�_�_�_�_oo %o7oIo[omoo�o�o �o�o�o�o�o!3 EWi{���� �����/�A�S� e�w���������я� ����+�=�O�a�s� ��������͟ߟ�� �'�9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� qE�_߿���'�9� K�]�oρϓϥϷ��� �������#�5�G�Y� k�}ߏߡ߳������� ����1�C�U�g�y� ������������	� �-�?�Q�c�u����� ����������) ;M_q���� ���%7I [m���������$PG�TRACELEN� sQ{A��� �&_UP ����H!�P 4!I !_�CFG �H%)2#!I �u$�@��/�,|@�*  ���%]"DEFSP/D �h,rA|@�� IN` TROL �h-�!8�%��!PE_CONF�Id �H%��H!u$4P�' LI�Da#�h-<PN6GR�P 1�+7� TP A>�ff��\!A�
=D�  DoZ� D\PA@�-` d�$�9�9C14P�;P�@�/�.�?G ´*CO�;B-@ TA4OO0OjOTO�O!�>�9S>��T�O�O�N�O =N�=m�h�O5_�O 2_k_V_�_z__�_�_ �_�_o�_�0z2c;o 
"ocooso�o�o �o�o�o�o�o)�&_J�n��z)��q
V7.10�beta1�& �A�k��qB
�Ӱ2�p?&ff^�q>.{�r��0�	����qB!��|�A{%�A��7�1�t �M�_�q�T��*�pu"�BȊ���͏ߏ�� α�O ��F�&��J�4�J:�KNOW_M  ��%p&P4SV ��9�;5 Po���h�;�&�8�Pq�u"�=O3Mx3�ɚ��0��2	�&BƠPV�ݯR��%�
Je�2�p@�0�� ,��(� ["LMRx3� ���F��Nc�E������{STx11 1�H)�4;5���;�> ݿ��2�%�7�I�{� m���ϣϵ������� 0��!�f�E�Wߜ�{��ߟ߾�2ɼ��ܿ G�<���y03����&ﾷ4C�U�g�yﾷ5�����ﾷA6��������7<�N�`�r���8�����������MAD%& �P&��OVLD  �H+֯����PARNUM  ̻�gy��SCH4	W R#
���	2#�UPD�eE5��_CMP_��% I �;0'p%MER_CHK[n#�"o�XjRS�@��P1_#MO6 ��_��տ_RES_GȰ�H+
:��?J/=/n/a/ �/�/�/�/�/�/�/?�?4?'?%��, '/Y?%B�v?�?�?# ��?�?�?#���?O O#;�3OROWO#�� rO�O�O#��O�O�O"V 1�̵�����P�|�THR_INR����z%dDVMASSQ_� ZeWMNP_�SM�ON_QUEUE� �̵�����*$NRU�N�V�X��SEND�Q��YEcXEo�UBE `|�_�SOPTIO�W���PPROGRAoM %�Z%�P�_��RTASK_�I6HnOCFG �ɶ_��o�`DAkTA����k��2��M_q��@ ������%�7�xI�[�~INFO���*}��T���ŏ׏ �����1�C�U�g� y���������ӟ����	��v����*| �E9�a� K_�a�8�i��]�ENB� l��	!��2����G�a2��l� X,	�	�=����'�@�"��$�����3TX�_EDIT ��oa�s��dWERFL"h7S���RCALL_CO�NF �l�F7%����ӿ�π
���KN�`?ڭ�����LDBD �1�P� /�)�C�￮���B6J` ������'�9�K�]� o߁ߓߥ߷��ߪ©� �ߡ��(�:�L�^�o� ����}������ ������,�>�P�b� t������������y� ��}�!3EW�� ~�������  2DVhz� ������// +/=/�d/���/�/ �/�/�/�/??*?<? N?`?r?��?��?�? ��?�?O#O�?JOy/ nO�O�O�O�O�O�O�O �O_"_4_F_X_3O|_ �?�_�_%O�_�_�_)O �_0o_OTofoxo�o�o �o�o�o�o�o, >ob�_�mo� ��o��Eo:�L� ^�p���������ʏ܏ � ��A�H�wl� S�������ß��}� +� �2�D�V�h�z��� ����¯ԯ���'�� .�]�R��s������� ۟пc����*�<� N�`�rτϖϨϺ��� ���߿�C�8��Y� k�}ߏ�����I����� ���"�4�F�X�j�|� �������������� �M�?�Q�c�u���� /���������, >Pbt����� ����3�%7I [��������� � //$/6/H/Z/l/ ~/�/��/��/�/ ??/?A?�/h?��/ �?�?�?�?�?�?
OO .O@OROdOvO�/�O�/ �O�O�/�O__'_�O N_}?r_�_�_�_�_�_ �_�_oo&o8oJo\o 7_�o�O�o�o)_�o�o �o-_�o4c_Xj| �������� �0�B�f��o��q� ��Ϗ���I >�P�b�t��������� Ο�����E��L� {�p�W�������ǯ�� �/�$�6�H�Z�l� ~�������ƿؿ��� +��2�a�V��wω� �ϭ�߯��g��
�� .�@�R�d�v߈ߚ߬� ����������G�<� ��]�o����Ϻ�M� ������&�8�J�\� n��������������� ����"Q�CUgy ���3����� 0BTfx�� ������/7)/ ;/M/_/��/���/ �/�/�/??(?:?L? ^?p?�?�?��?�/�? �?/O!O3OEO�?lO �/�?�O�O�O�O�O�O _ _2_D_V_h_z_�? �_�?�_�_O�_oo +o�_Ro�Ovo�o�o�o �o�o�o�o*< N`;o��_��-o ���1o�8�go\� n���������ȏڏ� ���"�4�F�!�j�� ��u����ӟ��� �M�B�T�f�x����� ����ү�����I� �P��t�[��������˿�$PRCAL�L_VER  �1�����WORK 2���:�
��\p����8ύ�( A� ��vψϚϬϾ����� ����*�<�N�`�r� �ߖߨߺ�������� �&�8�J�\�n��� ������������"� 4�F�X�1�Z�d���t� S����������� ,>Pbt��� ����(: L^p����� �� //$/6/H/Z/ l/~/�/�/�/�/�/�/ ��? ?2?D?V?h?z? �?�?�?�?�?�?�?
O O.O@OROdOvO�O�O �O�O�O�O�O__*_ <_N_`_r_�_�_�_�_��_�_�_oo&o߳G�ADJ ���/A�  Ve?��be��d��>bNS_C�FG �1���?�  BuzX�@��<@�0�?%DIAGX��o� 9��f�fveGRP� 2ڄgS` 	�HT�l�fn�{BP�`�@�`�2}*Fp/Hr **:QrASvs�d�"t X`Ȟ`1 An��{�m��c�x�qǜ���L�3�d�R�A�pT�4�.� @���d���������&� Џ"������<��� x�r����������ޟ �j��f�P�J�\�֯ ��ү����ȯB��>� (�"�4���X������� ���Ŀ� ���φ� 0ς�l�f�x��Ϝ��� ������^��Z�D�>� P���t��߰ߪ߼�6� ��2���(��L�� �������
����� � 8	 f�����<�����t$ ���������5GtgPR�EF ۄjs��s�
reIORIT�Y  p�Pcs���>aMPDSPON�  �y�b�UT��"swubODUCT_ID Ij�J�fOG�`_T�GL�Mf�HIB�IT_DO�-TOENT 1�Ij�* (!AF_I�NE� �!�tcp��!�ud��!iccm�w~�XY}c��d �s�)�a ^q>/P/s��8/ y/\%h/�/�/�/�/�/ �/�/#?
?G?Y?@?}?Hd?�?�?*�}c߄i¬b%a��?	Os�?+��<v^w/h|�?�ZOp���l�jA�b_,  �z bO@�O�O�O�xc�k�}�r>aPORT_WNUM�s���>a_CARTR�E)p#,tbSKS�TA�LSLGS6|�d��cs��Unothin�g�O�_�_�_Q�PT?EMP �Ii�_�=u�P_a_seibanRobo �oso�o�o�o�o�o�o N9r]� �������� 8�#�\�G���k�}��� ��ڏŏ���"��2� X�C�|�g�����ğ����ӟ��	�B��YVOERSI� �s�� disab�ledM�SAVE� ��
	26�70H774I�5�ϯ!JOѯ���C 	+��[�]�T�p�eq�������п޺A����	,��_W 1�d��P���$�Z�l�"�\ �URGE_ENB!E!WF��A���B�Wx��xA9ZW�RUP_DELA�Y �R^��R_?HOT %����IO9���R_NORMAL��(�}�L�SEMI\߂���Z_QSKIP8��WI�x3��/�*�<�N� ���m������ ������!�3�E��i� W�������w������� /��SAc� ��s��� �)O=s���/�$RA"��ۂL��D��_PARA�M��2��� @΁H@`�F�E2C��@�E�!C��FQB�BTIF�lTV\RCVTMO�UkWYU��D�CR8���� ���BL�B���-C�}?�0H�8"�8砊=���
S°���/�/]�� <
6b<�߈;܍�>u�.�>*��<ȃ��?{@�/V?g= �O�?�?�?�?�?�?�?�	OO-O?OQO�GRD�IO_TYPE � ?�G?]OEFP�OS1 1뛩�PxHOME�1�OB��%������(�>Ĳ��<ɛd���@���/_+_ *��O_u_`_�_ ��_X_�_|_�_o�_ ;o�__o�_�o�o0oBo |o�o�o�o%�oI �oF�>�b �����E�0�i� ���(���L���珂�����/�ʏS�e��E2 1����@���M�˟���m�S3 1턟�����`�K�|���S4 1���+�=�w�������S5 1ﮯ��ү����u���,�S6 1�C�U�g����
�C�>��S7 1�ؿ����6ϴϟ���V�S8 1�m�ϑ���I��4�m���SMASK 1�zO>#�߸ԋ�XNOwO��%�ޫA�MOTEL �K	�_ƹ����APL_RANG�O/Q�OWER �Y���["A��*S�YSTEM* V9.1060 ���11/14/2017 A �A0���n�RESTA�RT_T   �, $FLAG� $DSB_S�IGNAL $~��UP_CND����4�RS23�20��� � �$COMMENT� $DEV�ICEUSE��P�EE��$�ITY~��OPBITS���FLOWCONT{RO��TIMEg!���CUD�M��AU�XT����INTE�RFAC)�TATmUK���CH��� t $O�LD_/�C_SW� ��FREEF?ROMSIZ��_��ARGET_DI�R 	$UP?DT_MAP��R�TSK_ENB��EXP����! �F�AUL��EV���RV_DATA��  $$ E�a� �� 	$VA;LU9 	 ��_ z01A>"  �S� ���	� �$IT�P_6 $N;UM� OUP �?TOT_AXK��DSP�JOGL�Ir�FINE_P�C�j�OND|�$��UM{�K��_�MIR��P�T�N�APL��� _EX���������PG-BRKH����NC� IS �<  TsB^�P���D)�� BSO�C��N�DUM�MY162�SV�_CODE_OP�g�SFSPD_O�VRD]�LDl��OR�TP���LE�FU�� O�V�SF
*RUN�#��SF&&���U�FRA<*TOZ�L�CHDLY�RE�COV�#� WS0��|%� ROg��� _&    �@�@S5 NVER]T��OFS� CA ��FWD�x$���ENAB�TR����_FDO>MB_CM�� =B� BL_M���2$1���V�������3 |"G72AM�00��`5�"z?_M�60t�M{ tA�!T$SCA� �0D[�0�HBK�����1pE� �5IDX�2PPA�:�1�9D�5�5��1�#DVC_DBG��6A����7@�"��"NE1VJ�3NE3VF� /ATIO������U=C� �3j�AB� ��Y��� �$7�Y8��� _x���SUB�CPU��� SIN!_��3H4��1\73�H4��^$HW_�C1|Q�0<V��$AT��< �$U�NIThbP[PA�TTRI��oR� C�YCL�NECA��BFLTR_2_FI�1��C����{LP�CHK_��SCT�F_[WF1_e\�RwZFS��@2`RCHA�@�X/a?2i�.bRSD� ��x������0_T]8PR�O�@�#_�EMPER_� \TbP< �b��fDIAG~��RAILACDC�BMm LO{{!�M3�PS�h �0��E�3PR8@S�� I��qC*A�	�#�FUNC]��RINS_T����`�-t^�W�S_� ]�0Vs�п4VsWAR��2CBLCUR�kx�tA�{|Q�x|xD�AfWq�x�s�uLD@���1�s�`q�a��sTI�b	�< $CE_RIA��V��AF�@P��4�,� :�T2�`C��WB�11OIfP�&DF_�LETa� ��a�LM�B3FA� HRDYYO� RG�pHP`�����p��MULS�Ex���	W�`ap$�J�J�'�FAN_ALMLV����WRN�HAR�Dh���P��ap2��D�|@_s ��A�U��R!du�TO_SBR,Bq�� |�[P�,C5q��MPINFª qQ���q��RE	G�44V���"�#U�DAL_��FL=U]$M�p�P���	��0< ��4�8� � �� ���1g$YI����k|U��� �%�EG[Є�t�AR� �C�2�c���p2wAXE�ROB�
7RED�WR� Y_ӭ}SYV��[:��S��WRI� ��;PST���v�Z�w�nQ	��4�T�� �Bw�!F�5�c�0O�TO> � AR�Y�}��a�DH�F�I;|�$LIN]Kw�GTH����ST_<��!��6�NűXYZ��Ϻ7ݶ'OFF� ��Ĳ��%��B� "r"Ĉ!����#�FI�P<Ǆ�h��"r�_J�<����1I�U�_�8@�'�m`s�Ƃ��C��!DU�"��9�eTUR
�X��ŋ���1X��0��FLŰZ `�C����B�30�^�! 1> K� 	M���3Q�b	U�b	W��ORQf�\sP1ت�`8O�N�b����ّ��OVE��I�M���H���N� ��T��ָ��������� ��X�2'p�Q;�J��� � '�WB�������q�0N�q��ER�`qA	�b��#�c��A]�`P?�Nuzb���q�F�qAX�#<�q�@DQ ��	��a�ԁ�O�� m��ܰ����������1<������� !���1���A���Q��� a���q�����������ޢ�DEBU3S$�.q:��bR�"��AB��g�1���V�02R 
m_CJ���� �a�O��m��ܱ� ��������@���:�\E�#�LAB9���/P<CGRO�P��3��0B_�a��+�� 3�y�J~��zg��ANDP��@��Aɵ��g�� �1��ȱ�0�q��PȰNT�|#	 VEL�aC�!�a~&�SERVE	 Nc� $�ZpAk!!G PO�"3�0�w�N! 6"M�b�	�  $k"TREQ��
j#ޢt 
x'�:�2	�%��`_ � lpJ1�VERR_�82I�0 C�N�!TOQC�@�L��P���&z`GI%%�����4j#RE�p � ,E!�%� 
�G�RA11 23 dN2�3H,4� 7 C�$�Ѝb�j��*5OC�qt �  �+COU�NT?� IM��SFZN_CFG�s! 48Pۖ�RT���0S?AFP P�Q�x*1�1_� �� M�@�J��@?����@�%EFA'�N�5�)CX�ΠKK%I1I���J$��@ΡP�Bi HEL����2 5�k�B_BAS��RSSRږpȣS@����@17�@2�J3��J4�J5�J6�J7r�J87�AROOEИ0��ǰNLN���AqBV#�`�@ACK~KIN|0T�P�UI�8��!ajY_PU�S6��ROUX#P>pۘ�C�6"`�P��TPFWD_KAR�!�� REU$��P���qSpQUEڙz`�п��4�G�I���CŰ�c8 ͖űSEM�]ft���A!ASTYyT3SOH`]�DI�Q;pp�3%a��h�_TMMANRQ�fŰE�ND[�$KEY?SWITCH�S�Q�a.dHE��BEA�TMcPE��LEP�"SqfxU�SFLd��RS�dDO_HOeM8�O0�mPEF���PR(��2�,��UC�(pO��� 11OV_�M��3��IOCM���5g����FHKb� D±ܗ�0	U�"#bM|��T����FORC��WARؚ��"�COM�� G @\X�f�U2�EP��1*�/�,�3*�Q4y)2�0O�PL�y:2ۘUNLO�P��$x�EDL�  ��SNPX_A�S�2 0�AD�D�0�1$SIZ���$VA�5M_ULTIPZR���/�A� � �$�Y��\r=���S��39C� �FRI	F�B|0S`�`t��{NF�dODBU� ��P�K�U%�2�@c�� � ���"TqEӢҤ�SGL��	T���&�0��K�����STMT�ƓP�p��BW�Ж�SHsOWΕ�ABANڐTP�V��â�<ӢӴb�+0V��_G	B ��$PCS}0����FB�PR�SPR5`A�PT��8�D=�~B� ��!A00���3���=����G���Q���5��6���7��8��9��A��B��������B��F����^���1��U1��1ͩ1ک1�U1��1�1�1�U1(�15�1B�1O�U1\�2��2��2��U2��2ͩ2ک2穅2��2���.��2�(�25�2B�2O�2�\�;��Ȧ�������3�ͩ3ک3�3��3��3�3�3(�3�5�3B�3O�3\�4���4��4��4��4�ͩ4ک4�4��4��4�4�4(�4�5�4B�4O�4\�5���5��5��5��5�ͩ5ک5�5��5��5�5�5(�5�5�5B�5O�5\�6���6��6��6��6�ͩ6ک6�6��6��6�6�6(�6�5�6B�6O�6\�7���7��7��7��7�ͩ7ک7�7��7��7�7�7(�7*5�7B�7O�7\��r�VPpUq" z �B
7�F�>!��p}RaCM@@ "Mb R� �@$Q_�0R; �%�!�p�0#i YSL0?  � ��l��7;����Bp��;p�`�VA�LU�5�P�Vk�F��ID_LJ��H�I�I�r$FILcE_�S'$�T$]s쀠�SAp1 �h E@VE_B�LCKc`"��i(D_CPUy)��y)����3*/<$�p�RR � � PW��0LPS��!LAԑ�So1�#�!�$RUN_FLG5�$1�$@�`	5'1�$'1�%H�P��$I0�$$MC�TwBC2E ��� �`	0���Qy0.ped�4NscTDC	0�2�20@%��5�7THsF�3�]�6RLQyAESE�RVEfc�4sc�43�Aa1rP�0  �X -$ALEN`fc(Dsc@�PRA`L���W_y�#1A�$2bGMOq!��SF��PI�Pt !�IF�@�KDE�EB�LA3CE�rtCC��t p_MA���F�E�G��ATCV�LQ�GT �aZ0U&Zr��CY�TU$�CY�J�QU�MyT�P�J�W���E�Q�E'A2~`�|��Q�C��JK�VVK2��Q�q��QA�PJ&��Q�SJ�J�SJJ�SAAL��S`�S`f4e5�3�`N17\C`[�@
bL�@_@ba1�CF��! `] G�ROU����b^�N�x0C�`REQUsIR�2BpEBU��AzV$T�@2 ��a@�fa1��g4" �\�{APPR�`C�Lb
$OPEN�xCLOSJp"xSȸ56y�E
a1߆# �v�M�0�@BP��qt'_MG#!{pC��T p�x$��@�wBRK�y�NOLD�v��RT�MO_y3�w�}uuJ�p�tPd�@�S�@�S��@0c�@9c�@6�7�����qBg4$�# �bBB2�a��Qo�PATHk���z� ��GH����`#T;��SCAr�wrzqI�NBUC�@k�ڀC�t�UM�Yd@E  �P� !�1��P�@~�PAYLOA�w�J2LR_AN�1F�L� P�L�@�\���uR_F2LSHR�4��LOa�ف���������ACRL_@i!ׅʐӇ8�:bH��b$H�r��FL[EXs�a0Je6% P�bv?�?�?O�@}aJE& :'O9F�@����<O;a0�@EOWOiLF1��� �xO�O�O�O�O�O3�E�O�O __$_6_H_ Z_l_
�'�nW�S�T�@9ȍ_�_�_���ZTh��X���Uv�^��U �ű��_�_�_`ee�e0e9oKo]ooi_2J�d' �q0�o�o�o��0AT��axPE�L��Z2���hJ�`&v�`JE�pCTRӁ��TN7�־gHA_ND_VBb���U�( $|�F24�v�4�SWwbs��_v)� $$M n�ry[�q��q��Ͱ���r��A =�uv!D��~}A�|��zA�{AA�{���{� �zD�{�D�{P��G� ��S�T�w��y��N�xDY0p�v����^�@ ��������?��W^�ɠ���uP	���$�-��6�?�H�  u�U�* ��v�i���Cq��ASYM��t��`��)Tɍ��Ώ_ H0��߀��}�b���� �2�D�JK��p]�p}s|�)�_VIE���Cs�V_UN!I�3�ӈ�J�U� &������	$-&���xPΙ�pݟ%��L����i0H� �r+[�!'�rD	I�p�cO�$w� �ӧ, � �I�A  ����!�3 �/0�`0��  - �[ s�MEr�U�h#2}"
T� PT` Ћ�K1o`��&�B�P8k1_9Tata �$DUMMY1�A$PS_�RMFܠ  ���6kp7FLA�`YP���2�S3$GLB_T ���%�5K0r�X��'1. X�`�gU�SuT}Q�`SBRo �M21_V�bT$_SV_ERn�O5L!C9CCL�0!BA���O�"� GL�EW΂/ 4�`U1$YR�ZR�W�C�P��ro�A$0�A04dC]UjE0 |�N�@�f$GI+�}$jA q@dC�@��1 L�`�F4}$�F4E�FNEAR�l�N!�FYi�TAsNC!�1JOGР��p 2y`$J�OINT����bEMwSET�3  �GQE�E���S���D|�Ђ4� ��Ur�?��`LOC�K_FO��z�� B�GLV�GL�XT?EST_XMpwQ'EMPJP�b�R�2��P$Uj�iB��20�`�Ca1�Rv�Pa/#ACEq`�C#`_ $KARαM�#TPDRAm@@d7Q�VEC��Qf;PIU�a2aHE�PTO�OL�vcV�RENX`IS3b��b6$�N�ACH]P�`3�aQO��S3�43��@�SIr  @$�RAIL_BOX�E��F@ROBO��T?�FAHOWW�AR ��a�0�aROLM�2u~ѻd)r�Ѹ�`�W�O_F��!}F@HTML5�!"Ӂ�E�a�5C^0R[`O|�6CR۠LQ�PpSVOU_R7 	du@�U/
���ѣP_$PIP�VNj���b�b�a)�aspg�CORDED�P���p&PXT�p�A)� ���O
0 8 D �0OB&��ӨP1�� ��3�0 �4��SYS �ADR1� K0�TCH�� 9 M,|�EN�"0�A�Q�_�D����{��AV�WVA&1: �� F`jB�%PRE�V_RT3$E�DIT҆VSHW�R��F�j�~A��D50����$HEADEz "��UڃKE~A�0C�PSPD9�JMP�=�L�%��Rn��$Q;(�%���I�PS�ҍC?�NE`��5�T'ICK�l!M.�2P�a�HNA< @p*�����A�_GPЖ��f1�STY���aL�O�1�c�̒� =� t 
̀G��%�$���D=@S��!$���:1�5� �69PЖSQU:`֥<�2�TERCO0Azc@S��> �@�@��j���:�ma��OP0C3%�IZ�4�A�5�1PR��1�|��pPU���_DO�R��XS[PK�&A�XI�<saUR �Ћ����`��K�j���Y_m`]�ET^�P�R�9���F��A,����49�g`�0��SRR�?l�����£�ٵ��� ��ٵ��ٳ��ٳ��� ��$��4�1�K�a��1�o̟O�C��]�C�n�-?Qc_�SS}C�0 @ hF@cDSސAa�0SP� &K�AT"�����������2ADDRESz�cB݀SHIF��^�P_2CH0G��I�0���TU�0I���apCRCUSTOT�_�V�RI�"B~�P�X_�⣘ 
�Z
��qV�q�@C \r���x���ܼ�s�*�C�`󿢂����v?B*��TXSCREE"��D� 8�TINA\C�@}�D��_�_�� E Tr�<@�]� ;A@��+�\�+���ـRRO��(P03����4��UEh�F �Ț v��0S]A]�RS	M��!�U����&4�� S_�CT��D�W��r��_�C�R0�� �2Ex�UEGp�"LB���GMT@ %L!:�(@OMT��/BBL_�`W|0@�H ����O�A LE���`��
�RIGHBRD<ND��CKGR|0<�T�;8WIDT�H�c��2�1�1�a��IKpEY_���I��r[pp ��`�B�ACK���2�RA�.0FO�q�LAB�	�?(.0I�`�R�$UR�a� ��I_�40H�� J 8��!(P_!���50R�~@�R���h�1_��O�����KǐYG5 U�  `R�R#qLUM8`B��ERV�q�Io NE�L,0��GE��A}��*��LP���E���)�� ��0���`�5*�6�7�8���@C3�P>�6�a�Q�Ss�K�USR�jDM <r�40U��B���BFO���BP�RI��m�`N!� T�RIP�am�UWNDO�%N�@A��� #�
qX��R\�V� �O| �G �)�T<p����2OSS16Rb����#|a��PsO�C�ND2��v!�Q	U���QM?_?m��ߕ�#OFF�P��R�	@u3O�0 1�PF@�4�4QF@GUW�P�1r C��
G��SUB��U@��SR	TF0��Sǒ'QHpͣsOR�`PERAUҰQDTfI�����r��� T H*�SH�ADOW?��c�A_UNSCA_c�Ct��CDGD�a���V��VC�
`��U�# �b!�M�	d�N�a��c�C�p�EDRkIV�i�_Vِ�"T��pD]$MY_UBY\$T#�D3M���b�����X�a�R�P_�@���RL�B�M$��DEY���EX���aS�_�MUW�X�TI�US[�E`� h`��2� ����1G��PAC3IN��J�RG�*e�Ab�3Abj3Ab|��QR!E'��D1r�CAb�ppV ��TAREGGPP`�`�FR40�ppW�pY,�}0B	l�R�RE�SSW9`�_A:a�p�S�ODr!��A���cٲEM �U�)0�q�A�BHK�Xǐzv�б��`��CsEA��MwW�OR�e�eMRC]V��Y ��O �MCa�	�r�3�c�rREF���v�v~q �`����`� �z�q�z��q�{��v9_RCN{:�g{Y�SJ �WSSp����E��Z �񒠐 }��� XU��O�Uޗ~bߖS U�e��2V��~�@����W^�����Kn>�SUL X�3CO(�)Y�P�NT�Q��$��Q.�A.�i!.��L�SW��S0W�Ac�i!��D��[� ,^Ӕ�!н ^�CACH��LO�q�����PřB�l�~��C_LIMI�ӋFR�T7��t�$�HOwR��COMMS0�O &���0Ѱ���'�VP�b�`i�_Ӧs�Z%`n�n�WA��MP��F�AI�G?t��AyDépaIMRE���x�GP6��Pа�VASYNBUF�VVRTD�!�x�O�OL��D_�3=�W:j3P��ETU�SܐyQp�ECCUsh�VEM]`ԕ���VIRCá5��/�!�_DELAxc6�� �� �TAG1�R�QX#YZv�^��QW�a��d���T�@�RIM۱�4�����\�ҼLASj �q��_ܐ�>�I]�"ܑS堻�Nf�C�VLEXE���^��B�^��CFeL9 I�P�FI?��Ǥ@���T@s�� ������b_� ���z�:i#�Y ORD�!ȷ ��ӧ���U`���T�"��bvWOs _�@SFW �a  ���K.��P�URps�@SM�%yb�"G$ADJ1�f�U�����c�"�N�1LIN�30���|��d x�0MSPD$�B���J�	�p�rU��!��LNT:�B��M����*�NC��ACC�R'��SR�Q.� XVR�$e9����T_OVR���/ZABC=Ef�b���� 
��Z@�$gL�"�G$Lm�� ��_ZMPCF=Eht�����$��bQLNK�B
 ���P>Di �Ы3�Mp�CMC�M3`Cm�CART�_=�tPV� $J[�U�D^�a�r�`k��w���rUX � �UXE�Q�� �f���|�����������SP�Z��j P��m�4@��Y��D�0 kRѠ�!��HEIGH,cN�� ������P��l� � [�A��$�B�K�WgpK_SgHIF����RV�!F90�r���C� V�K� � b��5�I��S�D�TRAC�E� � ��PP�HERPm ,��8N`	��M�_DRY�%����k�%�,�|�[�`�B@ k���U �02i����P����! ���Gf�PR~�($(�#�2/D*R3�U/%&IcA_\�9�$$#��!_AIRPU�`  �  ����d�� �+��?�ISOLC  ��,�"�?����7;_$к�?���!H?774  f4�?��?�9[Z����#9x�[S232�� 1��C# L�TE�� PEND�A�`f4044D�f<]? M�aintenance ConsSB�1OSF"MO_DNo UseAM}OCO��O�O�O�O�O��2N�5��"31�%�1C�HP� �.,�	�	lQ7_!UDc1:�_9_&�AV��̻��%�"%�!SR  �+�`��_�PM�p�&�")`�.r�YV��!� 2��!� D�`P 	�/�o�Q�o�o�c ��o�g�o�o) M;]_q��� �����#�I�7� m�[��������ŏǏ ُ���3�!�W�E�{� i�������՟ß��� ��-�/�A�w�e��� �������ѯ��� =�+�a�O���s����� ��߿Ϳ��'��K��9�[ρ�oϥ���$�SAF_DO_PULS� �6Q���F��CA~нћ%6���R !�$!'A�,��0
@��]Q�4|A|E��b �oW�i�{ߍߟ߱� @���������/�*X+6S��2X�ъc�dX��b�:� @2;���������� }`���_	 ����T� ��2�D��V�c�T D�� c��������������� 
.@Rdv����_U�����	�
zC0B;�+o04p(e%�
�t��Di��0��/�  � �.60A/�'�њ �����//*/ </N/`/r/�/�/�/�/ �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4OFOXOjOoA���O�O�O�O�O �O�O_#_rOF�O_a_ s_�_�_�_�_�_�_�_�Q3_b0��}K� BoTofoxo�o�o�o�o �o�o�o,>P bt������ ���(�:�L�^�p� ��������ʏ܏� � �}O6�H�Z�l�~��� ����Ɵ؟C_��� � 2�D�V�h�z����_}[�S������	�����+���ί� ���$�5�G�Y�k� }�������ſ׿��� ��1�C�U�g�yϋ� �ϯ���������	�� -�?�Q�c�u߇ߙ�n��r�������� )�;�M�_�q����@�����������߸�E�O�����>�	1234�5678dh!?B!��,y���B�������� ��!3EK��n �������� "4FXj|� �]����
// ./@/R/d/v/�/�/�/ �/�/�/��?*?<? N?`?r?�?�?�?�?�? �?�?OO&O8O�/\O nO�O�O�O�O�O�O�O �O_"_4_F_X_j_|_ �_MO�_�_�_�_�_o o0oBoTofoxo�o�o �o�o�o�o�_, >Pbt���� �����(�:��o ^�p���������ʏ܏ � ��$�6�H�Z�l� ~���O���Ɵ؟��� � �2�D�V�h�z���@����¯ԯ��������?�Q�c��CH  Bp��_   ���2��]��} p�
����  	�p�2@ ������-����.����1��3 4 5 6-ρϓϥ� �����������#�5� G�Y�k�}ߏߡ߳���
T�(�������� *�<�N�`�r���� ����������&�8�J�\��� .�/�ʱ���<�� v�ʱ  �����]����ααt  �����]��$SC�R_GRP 1�!J!R�� �� �]�� ��	 /-�5F ?/�o�V]�R�n��s�����D� ��D�L��Q��	M-10iA�/12 1234�567890̰� 8̰MTC�3 *�
V0�3.01 Uu r�𼻲�|5�@$�$Qä?�C
x�	�����/�#/+$��H��5 �9$+!H����C}9�<��tC��X>���fB3CVB����Q¬PM���
�@�X����]B+G����Fr�~@?���C}2d�<?r�CϏ5 ׿�!��/�?f��/,;?vBǆ��W?U2�n4QA��}?  @0���5y?�7?��7Q2����?�:QF@ F�`�2 O�/$OO HO3OXO~OiO�O�O�O I=�1�2�O�O�O _TB� _�Of_Q_�_u_ �_�_�_�_�_o�_,o oPoB�`j��~g�o�i�
�o�o�c�1R#���o�0�4@�0���+w%%���kstA�yh�u�/�v �pQ��r�q  ����z�q�� +����a�s���o�����͏��ECLVLw  Ӂ�����r�L_DEFA�ULT�@ ������HOOTSTR��q��MIPOWERF��{��B�WFD�O� ��RV?ENT 1���:� L!DU�M_EIPӏ����j!AF_IN�E�ҟڔ!FT$���ȟ%�!X&A��L���q�!RPC_MAINr��T��`�����VIS䍯�����	�!TMP��PU ���d���U�!
PMON_�PROXYV���e D����o���f����!RDM_SR�V�gܿ9�!�RMtUϼ�h(υ�!%
��M����it����!RLSYNC�����8���!gROS��D��4ߞi�!
CE�?O�Mj߾�kXߵ�!	�~�CONS�߽�l���!~�WAS�RCϾ�m��M�!�~�USBN８n <��8���������� ���/���S��w�߇�RVICE_KL� ?%�� (%�SVCPRG1�~�����2������3�������4��5�>C��6fk��7@����F���9����P����3 ����[�����0 ���X������ �#/���K/���s/ ��!�/��I�/��q �/��?���;?�� �c?��/�?��9/�? ��a/�?��/O�/ ��������NO�O�� �O�O�O�O�O_�O'_ _K_]_H_�_l_�_�_ �_�_�_�_�_#ooGo 2okoVo�ozo�o�o�o �o�o�o1U@ g�v����� ��-��Q�<�u�`� ��������Ϗ�ޏ����_DEV ~���MC:��E�d1�GRP �2��5@��bx� 	� 
 ,���5@������ ��ʟ�����ܟ� � =�O�6�s�Z���~��� ͯ���د�'�����!�t�,��5@\��� �����ο��ǿ�� (��8�^�Eς�iϦϠ�ϟ���3�5@�5@ I��ϵ�>����F��� ��|߹ߠ�������� ��7�I�0�m�T������'���|���0��� ��%��I�0�m��f� ��������������! 3W��H�Hb� ������3 WiP�t��@���/���5@�5@Y��E/v// �/�/�/�/�/�/�/? �/(?N?5?r?Y?�?�? �?�?#/�?O�?&OO JO\OCO�OgO�O�O�O �O�O�O�O�O4__X_ ?_h_�_�?�_�_�_�_ �_o�_oBo)ofoMo �o�o�o�o�o�o�o�o >%�_t+� �������(� �L�3�\���i������ʏ܏Ï ��d ԿM6t6s�	� 9�o?b���@��ҹ��}?�P���_�*�>�����?��?���VrS�i#��@�zkE�¾}���W���
�����@«��xC,�E��g�M�HP`B��wA{9P@�r'���%�VIZPIX �1��$!�x%���.��qԈ�;����'}�Y �R>�������Q�������IAw�?����@a�4���n�¾|c��p��A,�����n]����C�&���4��?�FAY��@�ݝ���A"���%J?OGGING⟷��MQ6%�2Q�;�b�?�S�A���;z��@�fZ�il�������n-$@�z{@����A
#�A���9J��O����������bC�H�������&g��Bb~��vs��� ����P��ʟ����ɠ�����vv�n]_��e�,����>�\M���(��ￚ��1�����@�1�k[���9n?i��A�f�A�������C
����@�t%� ���AR��@۳���F�}A�Q�����\�Ǣ�%�_�>,xp>���}�"'��	�
�������@�;3��Ұ��l�GA�l\�9���!�mA9������s��LK�C
�<����������A����AJ��A(����3�e�w�!ߌ��S%�@9<�����G��k�:���=��?���=�2i���6ΒA����r���;���)��A��������A/�����l��z�C�	���>q![Aog�AvA}�)�Ag���w�� �Mn�ͥ�%�o���]>��Ы�=m���V��=*�?��Β������v��4>��G�A���F!����Fl�����¯�BZ�����������B�œ�AdLkA�ڛA���9ϸK���Ǡu�%����B/���v��/�:⠻��凉ā�@)���?���A������@�߯BB�Ye��d�������kE����Y�¬���C
&i����!?��A���-@�������~©�����N|���	M^�%����`f��ϜﾨW6�=#��v��.��	�h�AM�i�Z࿹��A�}| e��H���xu1A\���v��Ϙ8C��g����?����A_� AA��?6������~����Ǡa�������V߻��w��ÿ�"�/e���pǾ`�>A�6Z=�A�A�|qe���m?���2A$��Ȼ2$�ȿ�C7O,5��	>?��Aq��A@  ��?�D�א]o�TǠ@$%�=��qA�*�S�����9���$>�
��=�&��#x�@�"ѱ�@���H�W����A@�FA���]�(ͅ��y�C>�m��?��Ҿ���A@��A3��p�1A��h��="/aAm�I�,��Aڿ+\��+!�1�@��}�=����*��A%���@�TXA�������^�@�����?����=��C>c�����}��Ѕ1AK[��U��)�/X/�/gBp%�:&����6%�xu�~U"�|>w���>R�Z�3J��A��� H�@��V�8ӟ�e��(���E
�A<3������ȩ{Cc^�ν��?*���Az�B�z��eSAs�7��/�/�?ghd%���i"�k�o>���z?R�Bo?*������?�D3@�Y�L����@�l���_e��ϝ��vF@���3�2�_��?x)B���i����@��A�M@��[�K�AG~�:MAIN �?�O�0�%������{m�=�-��9:�=x ]���֓��@��@{\	A�`���#�A��i0O��n���0?a-��saµ�<C
��i�{-j@]�	>A��K���~AwƤ��y�O�Ox_�Ar���6#J�=�1�@H'Y@�ҏ��3��@����O��?�`�@�u5���C@���.���/��t��|�M����������ҟ�B�k�^=Q?��TA�̸@���A�`�mA�B�U_g_Lo ��P��6��־��t�@�wBA�Us�&S�@��]@�5�?k��)@1�����/�@�f�#�!|1N�m��Y���A	�+���Z�����B�y���@v'bqA�A�@����A<)oNo _a�s %�>�u�?�f±@���@��+˿]��@לȗi��c�2��@o"�����@�f��'@�8�y����k�{��"��Sۋ���KB��$�i������,��A���t������,AP*2��o"�3r�%��s��@���@���A*	@�����0ߍ�B�;|���Z@Cz�����:��Ag�݁~�C���̊A�k���^�ªM��C��i�� ���A���A|w-�?"`��T_��Ǐ^bvu�Y��C��oD�����:�� �ɿ��[/�<�=��� ��O�����'AW��~�X�'�0>��/��ʁ°�CB��X)=���@ ��A�i���="AC��F�e`*����ՆBU��Fb��<-f>�>���}�(���>���@�ɿ��@w������<�\��������޽�B�B�D=²�|�C g�N�>���ԙ�A�G�LA���A��i�y���p���D��u��k18����A�1��@����Ӱ�z�@�}ۿ����@st��٘��~��������A�β������4zB��N��4�䐺�A<��A��?�xA(|=�?�?�D��0L�I�mL�1=���=�d��G����W?�{�i�>������@PK_G�@֒�=�>�¶����	��A1#���u�v��#߬Cpf��������A���QA@����A�j02��V��XͽF�91����v����<��ɽ�l6�>� P��~�"����� ���7A��6��~�Yv�#�¿�3h����°(CӬ05=�?�����ABݝAv���æ�������W�[��,����cF��!@���"��ٖ�w?�c���R��A!���Q,^�@��[AT�z��~����y���ߤv�VW¸b�C$>L��eB�7>A��=�A7g*�	?K��l�M�;o~�� M]P����=��P@�r�@��?�ނ�ʁ�>�J$l?�Ơ@�`@�}o��#AY�H�_����v�@4����d�¹<��C�bu�7@2VA��m�!�@=�,����X���ߔ� ��e9u�?�zE=�|�=&kq����>�y�a���h��S�X@F0�a@��6��)ӟµ��W��uA����M��ƟP C�,����� �yA�.�?�Ư�����A�X�����h�W�]�s�a���8��+@M�@���a?oP���h�%�>=ք��@�fD3%A�$��A=�(jY��m�����@�	�����~¿���C0ǩ~���@7�A�L�A��@v��mwtq�k�<���h&]�a�@6��?�m����ϝ��@���*������@��@�9�.d�~��n��@���(E��̴C� CM������{A�3H�:�<�>Ac��>O:]�*S��@/ц?������@d|���?��@���=��v@�����#��~�q\����@��g���
�¿�/�B�H�?�'b���=�aA�z�E�2]A:0Єj��ID]�Z���@?�A��z���Fg@�=z�a.Kj?��P�@YN@�e?@i#����� ��e��I�@���:+D��Ð�B��>#C���㰰�i�@R&5��?�1A]�F����/O��@- �@Cl3?ѯ�=1�@+v�I�քeL�fA ��?@տ�!�5X�~����ݿ
@��E��?�;B��a�����rǭI��r���	�AY�Е/�/�?O�]�[���>|�1>iH��!��@�=^Q����@e�%�@�8�@_���bK��~�MP��^^�?-�n�E��[mB�+���������Aҩ���������A����i?�?`OO­�: ��@)�@_��2?�+@��i�7�Q�5����@h�0�Z�J���l@��P���so���N���� v¯�|�BO9���+��1��nlAZ��A��j���&�=ObO4_��n�1��bt��<|�*�36Q��2����~���0?�Z�}A!F=6Q!�A�AۑE�N�Nb����C��K���`Իª+|�C���;����@Z�;A�2�uAI�`�ԡc�4��_6_o�GR��պ�O�>�]�?����_I�!�S�����f��~�<� �D �A5�A��_N/��i߼��P�R�~�C�{Q�d��I��>Aɝ��A@���%��v���_
o�o��u����_�L�J��P��a<��>"@?	�Q��w�>�"A��@~��8����F�4�O����]=/?)��z�7�'µS�DBS�����@*��A���w��_�@��iA��ٹo�o�� MvK��I�;�?�/F?_��<����]@��A�Q�������{@c�9@�/����&��
Y��,��8��v��52��ߨC���= �������A��j�=t���W?D/AH:���섏�qzw��>�d�u?���?y��������=u��LQ��������@_<B@\��G?�;�=���n�����ߐ���-�y�CB�*Yѽ�����O�-A�$�Lk@dr'� �2�
m�R��v[��]��Z�@��?߬�2$R@%�G�-�x���g%2�%:��5!A1���<��A^-,=~�����Yݤ?l���APד­���C?.@ ������A�^����1�@�G����<5���,��k��]���@ ���@_Qx�*�h�?������ƭ�����@�ec5A?���V�=A�Y�=~���sI*>��ݧA�Q��Z:CC������A������ư@��x���<O���j��d]�d�=�n%=k��: ���@?���'ݰA�N�c�>f�@Ɣ��)����}���� AP�����A��KC��9��=}A��+A="c��?$�AUhE�W�\Կ+�e���2���>���?�U���&i���x���*p@!�����m1�(�����TAAW�Z���(�������e��¨�χC���b�V����ҖB����AM�p�8���ÿ��粩��5b>��?A�2i?,��������L@� �f�����t]1�~C�/����Q���JYϟ`>����&.B��AS�-��ϔ�y���n���=���<�c�v<�:�'}1�=$D�����T?3J�:Ձ>����m����"���I@���|52���C����P��n�A���A9P�=��t�AP��yݯ�P� (M�By6T�r5��T�3������):� ����@��\��yS`��AV:��@��dZ�k.��D�B.�ZA��h{���¿�Z�B���>@�N��+�������A�_��(��@뢠Y�k�$���GA��>|�c?�����Ϗ"��N���y�����@�w�����A<Iq����2�mTO52��_C);�Ο�![�� �����A@k��}���-������_u���v�o�<͚�%?���?�b��@CH��z�� ��T�W�Hb�o@�9��2 �w�A$:�=~�H�X�(�$���kK�m�����B�jm.�R�0�7��B�A�AQ1�����B���	SCAN_SL�OT���M_z�;MV�#@0�@I6�>�����>�4?�r��@8���0���@����p��@�t]�-��n�=���=��[�ו#?����y��@�c�G��~ �+m�B�	QyAwg*�6��Ac�	���� � QMU���RU@%6�@�p>�=���������n@�:R��R`@}�����*@���"A*�
=~Bw����r������>	}/�~A��BT�޾�$��mB�zA������b��GC}�t/�}�v��v� �?���#5bTɿ��Ž�D�v?���@N ?������3�A����Z�4��������2$��SBZ��=�NC�?�-�jA!@Ư�A?e���_Q/c/�H?��MU��o���@B�����ưҿ�Jd��^��?��Є�{���<�Y���AKg=~F�A�������r����]� �BF� .>�	>�@��BU���[�@�1�W %?7?O��{'�v��k?�ߑ&@�zr?���I@K����7�����f@u�5U��oTX��ZT�=~� ������wy��aY#y���?'��M��9>KBÞA�*��J^A��~�
CHECKO��O1@@MU��O�<=<C@]o��5b����(���m^����*��@��}=^aߔ�Ah���<���'��(����V������]���0��#��1A�ʂ�@'����+��O�O�_Q~-�v����@C��@r�b0�D�6?�?�?%͍������7@h�.�A˞�f��b�=}��A�k�$Q�7�/7z��&�e�"��n?�<�bA���
��.A�#IA��(�[BLABE�L�_�j	�P�	U��9���Y��:��_-��^��aa�����9q�@�y@����@�3�A���=~�iw@�k�������F��«:$��[,�������[A] j������q���/�$;�ognsMa0�/	U����<��H1=h�>����=֝۾=���@&�����|O�������|A�Id�i��� ����-�������><�y��Іs������  'B�p�@��\Av?��|�?�_�@��a<�	U��O�L��M�/o;~�m/xϿ����{\�	AU[��e�?@�1AP+��a��`������@>���r���H��'��ޥ��@_��BA�Z)A���A���������I[� U����v�����]��%E>h�����bW?i)�����˿A?��Y������	�a���@����A���>9.��?v����]�^`�@���A��-�Ak��>��A(|�*�_��Fa�Tj	Ps�B�P��?�m�?�uG�=��?Q��@��d��v�@������Yv��G�la��V�����h�U�'������Äć�N�����1�A�o@�A_��AK��AǾ�LI'GHT���#���#�۰M?�dD?��D�=6��??%"�@���
aE�r�9�~����Eu ��$���7v��U�4����Å,/�N�������A�AbcXAO[��AzIA��DEMؠ�qTl��U��?�ų?rY��;�*�?�@zC��|=��`�@[��I�ͨe����J�{֠Z���������u�U����%	���Å����B� ��yA��?�w�`A&�y6�VIZPIX���f���mզ���?��4?���;��&?8
��@�v�1q�߿�,^@FQ5���Ō��V|���b��t���U�'��<���>Å�����(I��O��A��@��A��xA�ڡ�A�S�8�w�s�`���ҡ�1=�/��=����~�ܿ����N���`>�az{>��k��<Aa2���~��(�����`�׹�����¾{��UC��ǯ�A��@A����al���3ş�ן��Pm�4	P�=y��������?��d?[7.�nvD��@��AX�A�Q��ec5����[AQ��~M�,�sC����(�A���e���Y��).���0@�qA�R�A���������������P�
v�=����D߿b	:v0�����<��Z]��������hA-��%AEw@V��=@�n�~���F�������?��K¥���CMb�Ng�M@=�A������"c��?�i�Tp!�'�ܴ�'�
x�	U=������7��+c�f?�7�x1)����N A*�*=(���@[���H4��A��|��������9���¬E�C ��?ڀ?� Au���A>��ƒ}�A�}l�����z�	U@,��@�+@ 7y<��¾;L?��F��.=ք�U��U����J@��N��"���������G�A�6��)N���3C���N�0Y��i�A�W���]j�AQ��ew\ )� ����?`l@���ǡ"�J濲���>b���"�@�6�b~ͩA>��	�~�\���o����
c���«7�C��i�>���m�PA�KE�����Aڛ����9K0/ � ��	U:j0?l-�@��En�'}?��L��Ch�N�rA���1A����z�OA3U���\���J7��W�g�vO�­��C˦�� ��aB�A������oA7��`�x��/�/=(�զʹ����s7�-�q�:n����?�2�f�;3��	��A�(�@e�w��Hz�����!� YA!�I��%f��ȓ#�C�H���@2VA��R�A����B��AB�d�/�?  _M
|	P2����R >���?v��Q�>�삾�fڱB��?�d�7���mA��S@��mA�0�t�/-Z������©W����¨=�C��8�H�!�=���B�>����9P�>�V��Çy�?�?�OC!|���fj�?�@�@�j#��`?������QE�hw0��aKj-A���jA8�P��~�}��S���A ���D���{�Ca���Z�;����A�O��ư�@Y���r��X�O�O�_ $�0�Y��Wp�+'�����<cR=�(�Ͽ�z�?2�i��~ A�#���#���f�A,1��~�>}��͔�A5U��9U����Cxѕ�*�?4��A�1A�~� !�_�['��i_NoVdM
~0���>ǐi?�7�$B����n� ��"�����@mL%@������C�A-��9O`Ŀ�S �@S߾�$»�C�n�?���
%������F��f$�$1oCo(C =��Y�Q��nP��S*Q<uZX�=<������VrS	A�X���v��t�]A1id?�Q���ЭA3�w��P� ����C�(�}� ���>�![AN���A��A4���k����g`Humj���?�O���>�?���W�~�P�����@x��A
4,A�AR^��ʓu������OA���p�­�mC�^���� A�N��w�vs����4�z��ʏ5wH}�9��ǿh;7�hb�|�`xȼz��
?�^U�
 ����ٱA5D��@��q�(����ow�?�yA�/���.S'�?�QCez���p����AgW�C��@��%/AW}�*���������զ������<��ý�^ �.k(?>�)�Oja�� A���ѿ�d���O��������X�A/�_�������C+�CU�z٢�����q�pb+�A=�"c@�e�A�������x���n��E>�"9>7>� F:^ ;���=��^��^᭔%@Q,^�?���@�'��E/����=��?�8A0�������l6�C��E�`��U�A�m�@��ư�L�A��L�U�g�L�oq����VE����9fн>�4�="����z ����7Ar/@���@{�e����ٯN�@ ��A09�l����nC�l�JP�A��z�@Bݝ���A/ώ)�;� � �(Mw1�E�w��Ͼ%YD�*�E<!�<׿LF��-������������m1����A-�J�����6�����A6�0��#���C��	o�}��߈A�g*)bo�0�
	���	�x��E�2�g�?���B�]��>����� H@p��@�� ����A4�Xm��Q���K9�@�a���¸�q�C������A�����IAF�}�iͰ������݇y�E9�R!y��@����}����RIޱ~`�>��@���A�%�#��U�R����h��d�d�$s�­A�C���m�=�pIRɝ����H�A����h�>�߷ߜ������~^���^� ���[?�!��}޽ք�]z�EA'4�@��@mD+�x�|)�R����`��: ���/®��M�7��>�}=�q�ϝ���0�;A�y﬋�p� ��J��}]G��哹21�e�?�ѹ}��}����A�)gmA �?@<��	�_��a��R|�@�6�3®�e�C����ݿ	>>��!=��������A-���M�_�D��>��u�G@O�l}�=a�;K��}�Dp�X@�u5A0���d0AL��]��ͦ��:�[�'����­��Cié������[A�������A1?|"���!3��C�V=c��������~<���=E�d�� ��^�m������}����A5��~��.�XlgA�1-w�yi�pq߀Cz������=�Au��A�?W�A"�MY_���c@��Z�ߘ�1v���F?Qu�Q�~p��k�)A�?�!�@�����'�~�9M�y��r@��߾���L¾-C���-��p?]	>A��eSAH���6������/�i�9�!��.=ｼ���;D8ߍ��D�^[��I����A P��@���@rlߛAD%�~�^����\A6���(ͅ��*��C�5^l�T@FnMR����On�߫/�?��e9��?�����>��g�<��cR<� ]�+(�X�?: �����.��[��A�IP���8w���~KA6E6��2����nC�� ��� ?����AtC�A
�{�@F���_Tq?��?hO�h8�2�q;�NO�?�.�@��Ҵ<��@,��r����h����?�����,^�:��A5�BM/�o�������+C���¥���C���ARb�F���TB��U�A��:��VD�EOWO<_�P�h6�Fb�?f�$(@���;��}E?�F�����y-޶Β��N/?�\	<���!�A���n��@���f�������¥��gC��ݞ��C��2��B��h����Bz?14���<_+_�o %}@R]	���`��DI�<P�ϝ�~yW@A�|-�j��"���.h@����o�\ pw@���A��������?��#C�p:���F���A�`��A��g���AP*2�Z�JOGGING�o�nMpc�E:�w��?��@��S�<���@v�I�,/-��2��~�@�T�W?AZ}����A!5T������Ӭ+����p��+�¥���C��ݞ�������B�����-z�<�a[�_�_�+s8�ݾ��vwx鱾�?5�>�?�ݝ�Q�m�%:�@mL%�@����:yt�E������Σ����}¿���C������!�A�9��l��A�b�JA�+w�o�o���`4�պ΋@ŗ�?�U-�6����*j=�f��-�����
�@R�Z������_ qo�ؿ���rA/�־��=���C�Ĩ�@�=�����A�A���&�*t�AǠ>���`� !�M6�ٽ�`�����M��>v�뾯A!AB =���>@��R����Ďº*<�E���l�����²XvBM�k}��?��0�I�`�"�RW�i�{�4���6:�?�VYy@�j�����?������-ޖ���t@������MIsA�+�x�$��������u���.�«!5C�
	�
 � ��A���?�v�@�TY�^4�p=�O����6a1�K5?������f�<jP=�߲��/vQ/����QAt]����V�}ŒA)�r<����,�����wA3�L������ʰ�C�x��NR�0?���Ab+�A���A?C�]c�F���ܿ Q��$SERV_M?AIL  �ѽ��������OUT�PUT ����@��RV 28���� (a���0�޿h���SAV�E!��TOP10� 2A� d ��  �UR  ���I��]�6 %*�� ���sZ��� ��I��%�7�I� [�m�ߑߣߵ����� �����!�3�E�W�i� {������������ ��/�A�S�e�w���`����������YP����FZN_CFGw ����V�u���GRP 2��� ,B �PE qD;� B}P�  B4hÿRB21t�H7ELL�����ƈT�U�h��lRSR���	� -Q<u`r� �����/)/;.+�_��I�%;/i/P{/I"�,0�� �/��"� ހ'Q"��d��,�-��pHK 1~ �/ ?*? $?N?w?r?�?�?�?�? �?�?OOO&OOOJO�\OnOjOMM �~�OoFTOV_ENB��I����"�OW_REG_U�I�O�IMIOFWDL�@�NHR/WAIT�B�)�;V��FH�8YTI�M�E��r_VA���I_Q_UNIT��C�V��LC�@TR�Y�G���@MO�N_ALIAS k?e�IP�heH� o1oCoUogoqfo�o �o�o�ouo�o $ 6�oZl~��M ������2�D� V�h��y�����ԏ ���
��.�@��d� v�������W�П��� ��ß<�N�`�r�� ������̯ޯ���� &�8�J���n������� ��a�ڿ���ϻ�!� F�X�j�|�'Ϡϲ��� ���ϓ���0�B�T� ��xߊߜ߮���k��� ������>�P�b�t� ��1���������� �(�:�L�^�	����� ����c����� $ ��HZl~�;� ����� 2D Vh����m ��
//./�R/d/ v/�/�/E/�/�/�/�/ ?�/*?<?N?`??q? �?�?�?�?w?�?OO &O8O�?\OnO�O�O�O OO�O�O�O�O_�O4_ F_X_j__�_�_�_�_ �_�_�_oo0oBoIc��$SMON_D�EFPROG �&���la� &*SY�STEM*Io�g�@�P[dRECA�LL ?}li ( �}�_�o�o�o 2 �oWi{ ���D���� �/��S�e�w����� ��@�я�����+� ��O�a�s�������<� ͟ߟ���'���K� ]�o�������8�ɯۯ ����#���4�Y�k� }�������F�׿��� ��1�ĿU�g�yϋ� �ϯ�B�������	�� -���Q�c�u߇ߙ߫� >���������)�� M�_�q����:��� ������%���I�[� m������6������� ��!3��Wi{ ���D��� /�Sew�� �@���//+/ �O/a/s/�/�/�/</ �/�/�/??'?�/K? ]?o?�?�?�?8?�?�? �?�?O#O�?4OYOkO }O�O�O�OFO�O�O�O __1_�OU_g_y_�_ �_�_B_�_�_�_	oo -o�_Qocouo�o�o�o >o�o�o�o)�o M_q���:� ����%��I�[� m������6���ُ� ���!�3�ƏW�i�{� ������D�՟���� �/�S�e�w��������@��$SNPX�_ASG 2����ӡ_�  0A�%G����A�?�ĦPAR�AM ӥ^ݡ �	�P��eA���O��Ơ�OFT_KB_CFG  @�٥ã�OPIN_SIMW  ӫJ����ȿҳƠRVNO�RDY_DO  �T�|��QST_P_DSB��J�|(ϻ�SR ө� � & C�HECK_SLOT �E4���u�Ԡ�ƠTOP_ON_�ERR�Ģ��PT�N ӥ����A��RING�_PRM���VC�NT_GP 2tӥL��x 	$π#�A��J�5�n߿�V}D��RP 1#�M�_�ϱQߩ߻��� ������'�9�K�]� o����������� ���#�5�G�Y�k�}� �������������� 1Cjgy�� �����	0- ?Qcu���� ���//)/;/M/ _/q/�/�/�/�/�/�/ �/??%?7?I?[?�? ?�?�?�?�?�?�?�? O!OHOEOWOiO{O�O �O�O�O�O�O___ /_A_S_e_w_�_�_�_ �_�_�_�_oo+o=o Ooaoso�o�o�o�o�o �o�o'9`] o������� �&�#�5�G�Y�k�}����PRG_COU�NTq���¢�ENB�Ϥ�M΃s�ۏ_UPD 1N�T  
��A�%� 7�I�r�m�������� ǟٟ����!�J�E� W�i���������گկ ���"��/�A�j�e� w���������ѿ���� ��B�=�O�aϊυ� �ϩ����������� '�9�b�]�o߁ߪߥ� �����������:�5� G�Y��}������� �������1�Z�U� g�y������������� ��	2-?Qzu��������_I?NFO 1���� ���?�
��?��&@	���������@�ℌD��@C@B�C����| CR��@=?�d?�ц]@�����>(�	��?����q-���BO�o����	2z	���Q��YSDOEBUG����� �d���SP_PA�SS��B?�L�OG ���  � !?��� �  �����UD1:�\$�"_MPC�/ @$C"�/:,�J(2V/h"SAV �)($�*�J(SV�TEM�_TIME 1�'� 0 ۰y����  ���'.���7SKMEM  ����+  �  � %�/�?�?��X|��[BwF : d"�5�к?O pH�D0� d0OAM� qG"�WE���!�AG@BzO�O�O  �MgK�E� ��OjJ�O_U�V� �OH_Z_l_~_�_�_D�_�_U�_�_��e�_ o/oAoSoeowo�o�o �o�o�o�o�o+�=Oas�T1S�VGUNS���'�����pASK_?OPTION���t���q_DI��Ϗ�uBC2_GR/P 2��52��pC' C��||BC?CFG !�{�-1�"�/U�`s�? ������ݏȏ��%� �I�4�F��j����� ǟ���֟��!��E� 0�i�T���x���������֬�ׯ8�J� ů'���k�����ȿֺ 쿾p"���:� (�^�Lς�pϒϔϦ� ���� ���$��H�6� X�~�lߢߐ��ߴ��� �������D�*��X� j����*������ ���*�<�N��r�`� �������������� 8&\J�n� ������" 24F|j�V� ���/�0//@/ f/T/�/�/�/|/�/�/ �/�/??*?,?>?t? b?�?�?�?�?�?�?�? OO:O(O^OLO�OpO �O�O�O�O�O _�_ *_H_Z_l_�O�_~_�_ �_�_�_�_o�_2o o VoDozoho�o�o�o�o �o�o�o
@.P vd������ ���<�*�`�_x� ������̏J���ޏ � &��J�\�n�<����� ����ڟȟ����4� "�X�F�|�j������� ֯į�����B�0� R�T�f�������v�ؿ ���,Ϫ�P�>�`� ��tϪϼ��Ϝ����� ��:�(�J�L�^ߔ� �߸ߦ����� ���� 6�$�Z�H�~�l��� ��������� �ֿ8� J�h�z���
������� ����
.��R@ vd������ �<*`Np ������/� //&/\/J/�/6��/ �/�/�/�/j/?�/ ?�F?4?j?T6�0�$T�BCSG_GRP� 2"T5��  ��1 
? ?�  �?�? �?�?�?O�?	OCO-O�gOyK�2�3$�<d�, ��A?�1	� HCA�wE>w����B���wE?CS�C�2�O��H�JuR�M*��O6]B�yH�0TR3[33wEBl�@6_~]A�yH]Q]P�I�Q�C\~_�_yH���V�_o�Y yO,i aC�oVm@UQPMih |e�oZolo�o�o�o�o�.{x�a�	�V3.00�2	�mtc3.s	*�jpbt�2y8v�QY�ٚ�0!` Hy ��p�}�  a@���͂��u�1J2ʓ3%�=��CFoG 'T5�1Y �00��Z��r90�������� ��]0��ߏʏ��'� �K�6�o�Z�l����� ɟ���؟���!�G� 2�k�V���z�����ׯ ¯ԯ���1��U�g� �2� r�����@�ɿ�� ٿ���#��G�2�k� }Ϗϡ�\��ϰ����� ��߈1t?D�P?T�V� hߞߌ��߰�����
� ���@�.�d�R��v� ����������*� �N�<�r�`������� �������/,�� Ln\����� ��"4�DF X�|����� /�0//@/B/T/�/ x/�/�/�/�/�/�/? ,??P?>?t?b?�?�? �?�?�?�?�?OO:O (O^OLOnO�O>�O�O �OzO _�O__$_Z_ H_~_l_�_�_�_�_�_ �_�_ oo0oVohozo 4o�o�o�o�o�o�o�o 
,.@vd� �������� <�*�`�N���r����� ��ޏ̏���&�8��O P�b� ������ȟ�� �ڟ�����F�X�j� (�z�����į����� ��دB�0�f�T�v� ���������ҿ��� ��,�b�Pφ�tϪ� ���ϼ������(�� L�:�p�^߀߂ߔ��� D�������6�$�F� l�Z��~������� �����2� �V�D�f� ������j�|�����
 ��.R@b�v ������ N<r`��� ����//8/&/ \/n/�/�/�T/�/ �/�/�/"??2?X?F? |?�?�?^?p?�?�?�? �?O0OBOTOOxOfO �O�O�O�O�O�O�O_ _>_,_N_t_b_�_�_ �_�_�_�_�_�_o:o (o^oLo�opo�o�o�o �o�o z/�/*<�o Zl����� �� �2�D��h�V� x�z���ԏ����� �
�@�.�d�R�t�v� �������П���*� �:�`�N���r����� ̯��ܯޯ�&��J� 8�n�\�����N��ο ࿊����4�"�D�F� Xώ�|ϲ������Ϧ�����0��T�>�  9z�~� ~֒��~��$TBJOP_GRP 2(F���  �?�~�	�ұ�*����N��_xJ�Ќ���  �<� ���~� �@z���	 �CA��.��SC���_~�����>�f=fR�?��N�`��=#B�CS��?�l��z�?���C4  B��D���.�@�?
=�q��333����;W��h��$�l����R��Ҙ�9�����N�C�  D\"���!G�r�Ll��r���;L��Bl�  @fff@�>l����C���L.���A���Z������#���
;1U�x��@��p��?�33C���z ��Y����`���ޠ;xCs2)���@;�@VffB�f �zH�w�R".{�0:�t-�@	
� 0��p���t�� ��������/ ��$/>/(/6/d/�/ p/*/�/�/�/�/�/%?���~�bzиJ�	�V3.0[��omtc3��*p0���y�~?�7 E�o�E��E���E�F���F!�F�8��FT�F�qe\F�NaF����F�^lF����F�:
F��)F��3G��G��G��G,I�1�CH`�C�dT�DU�?D���D��DE(!/�E\�E���E�h�E�M�E��sF`�F+'\FD���F`=F}'��F��F�[
�F���F��M�;��
;Q��<.zГ� f�*���nO�B~��C?������O��ESTPARS  r���Ч�HR�@ABL�E 1+�� $�@~��H�G �yI
�G�H�H}ׅ��G	�H
�H�HU~��H�H�H7 �D'RDI�O��_$_ 6_H_Z_lU�TO�_�[@�_
oo.o@n�BS�_�� �Z%7I [m����� ���!�3�E�W��� �`�o��W���o�o�o �oc_u_�_�_�_�X�B~~�NUM  Fի��
��� �P7 �B_CFG �,g��"�@��IMEBF_TT�A0����@��VE#��Q�������R 1-�[ 8{?~�dy�� IУ�  � �(�:�L�^�p����� ����ʯܯ� ��$� 6�H���l�~�ǿ����ʿؿ���A���&���MDH�Z���ϐ��� V_I���Ϥ�GINT��ߤ�TF�8�J� B��d�vߪ��_TC�ߪߤ�	$0�@����N�RQ��R�_a�֖@���@MI_CHAN��� �� ��DBGL�VL�����A��E�THERAD ?��E����@0���:e��4:41:8b:b9 ���a+��`��c��RO�UTӐ!ej!�8�V��I��SNMA�SK������255.��\3�������\3�@OOLOFS�_DI�@P��O�RQCTRL !.�Lc�O4T#X j|������ �0BTfx��"����CPE?_DETAI�����PGL_CONF�IG 4g�w����/cell/�$CID$/grp1�I/[/m//�/Gc���/�/�/�/? ?�/:?L?^?p?�?�? #?�?�?�?�? OO�? �?HOZOlO~O�O�O1O �O�O�O�O_ _�OD_ V_h_z_�_�_-_?_�_@�_�_
oo.o��}�_ dovo�o�o�o�o,���o�m��_-?Q cu�_����� ���)�;�M�_�q� �������ˏݏ�� ��%�7�I�[�m��� ����ǟٟ������ 3�E�W�i�{������ ïկ������/�A� S�e�w�����*���ѿ ����Ϩ�=�O�a� sυϗ�&ϻ����������'�" �U�ser View� 7)}}1234?567890X�j� |ߎߠ߲ߺ�C�#����>�2Kٷ��.�@�R�d�v�����E�3 ������������}�?���4��x������� ����1�����5g�, >Pbt������6��(:�[��7����@���M/��8� H/Z/l/~/�/�//�/��" lCameraI�?/?@?,?>?P?b?@bE�/ �?�?�>V��?�?�? OO$O	  �&���/ tO�O�O�O�O�Ou?�O __aO:_L_^_p_�_�_�/��&��+_�_�_ oo(o:o�O^opo�o �_�o�o�o�o�o �_ �Wf��oL^p�� �Mo���9�$� 6�H�Z�l��W@K� ��̏ޏ�����8� J�\�����������ȟ ڟ���%�	o�$�6�H� Z�l�~�%�����Ư� ���� �2�D�럹W �ۯ������ƿؿ� ��� �2�}�V�h�z� �Ϟϰ�W��W6)G��� � �2�D�V���zߌ� ������������
������9��]�o��� ���^����������5�G�Y�k�}���*	�%0�������  $��HZl��� ��������� �+ �CUgy��D ���0	//-/?/ Q/c/
�%WK��/�/ �/�/�/	?�-???Q? �/u?�?�?�?�?�?v/ ���[f?O-O?OQOcO uO?�O�O�OO�O�O __)_;_�?�5/{�O �_�_�_�_�_�_�Oo o)ot_Mo_oqo�o�o �oN_�5��>o�o );M�_q���o �������o�5 ��_�q��������� `ݏ��L�%�7�I��[�m��&�   *�����ҟ������,�>�P�b�t�   }��?fffBhP���&�C"���-�QC���?���SB?u�A��h�>���g�D��D,g��� r������0�B�T� f�x���������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ���߸������ߜ�  }
&�(  袐( 	 ��,�� P�>�t�b�����������:� ��� �Ώ����� ���������!(� n�K]o����� ���4#5| Yk}����� ��B/1/C/U/g/ y/���/�/�//�/ 	??-???Q?�/u?�? �?�/�?�?�?�?OO ^?;OMO_O�?�O�O�O �O�O�O$O6O_%_7_ ~O[_m__�_�_�_�O �_�_�_D_!o3oEoWo io{o�_�o�o�o
o�o �o/A�o�ow ���o����� �`=�O�a������ ����͏ߏ&���'� n�K�]�o�������� ��۟���F�#�5�G� Y�k�}�ğ����ů� �����1�C���g� y���ү����ӿ���8	�P�0�@ +�8��J�\�+�2�����#frh:\tp�gl\robots\m10ia��_12.xml� ����������&�8�J�\�n���nߓߥ� �����������#�5� G�Y�p�j������ ��������1�C�U� l�f������������� ��	-?Qh�b ������� );Md^�� �����//%/ 7/I/`Z//�/�/�/ �/�/�/�/?!?3?E? \/V?{?�?�?�?�?�? �?�?OO/OAOSNuȝ�� 2π�<�< ~� ?� SK�OSO�O�O�O�O�O _�O,_J_0_B_d_�_ x_�_�_�_�_�_�_�_�oFoT��$TPG�L_OUTPUT� 7^�^� v@�e�o�o�o �o�o�o'9K ]o����������#�5��ev@��K`2345678901Z�l�~����� ����T�W������ +�=�ՏA�s���������S�}ş����#� 5�͟ߟk�}������� ů]�ӯ����1�C� ۯQ�y���������Y� k���	��-�?�Q�� _χϙϫϽ���g��� ��)�;�M����σ� �ߧ߹�����u���� %�7�I�[���i��� ������q���!�3� E�W�i��w������� �������/ASe��Va}qA������@xO*<�~J ( 	  ?�q_����� ���/7/%/[/I/ /m/�/�/�/�/�/�/ �/!??E?3?U?W?i?�?�?�?M��t@�F�? �?M�?1OCOOgOyO G��?�O�OVO�O�O�O �O(_:_�O>_p_
_\_ �_�_�_�_�_L_�_$o �_oZoloFo�o�o o �o�o�o�o �o, V�o�o��8�� ��
��z@�R�� >���b�t���Џ.�؏ ����<�N�(�r��� �l���̟f���ܟ 
�8��� �n������ �������J�\�"�4� ί@�j�D�V������ ��迂�Կ�0�
�T� f�ĿNϜ�6ψ����� ����x��P�b��� �ߘ�rߤ���,�>�� ���L�&�8��� �߸���d�� �����6�H��2)�u���$TPOFF_L�IM �0 �1����N_SV���  ��P_MON 8�5S��  2���STRTCHK �9�5��d���VTCOMPAT���D��VWVAR �:��g�� � �������_DEFPRO�G %		%
�CHECK_SLOT RAME����_DISPLA�Y��	�INST�_MSK  � �
INUSE9R:�LCKC
�QUICKMEN�g�SCRE���5Etps�c�C����_�ST8
��RAC�E_CFG ;���g��	�
�?�(HNL 2!<�
�0&!n �Z/ l/~/�/�/�/�/�/�*�%ITEM 2=�F+ �%$12�34567890<-??5  =<7?]?<o?w3  !}?�;� A?�?�+?�?O? O!O�?7O�?�?�O�? �OO�O�O[OKO]OoO �O�O_�Oc_�_�_�O �_#_5_G_�_k_o=o Oo�_[o�_�_�_o�o 1o�ogo�o�of �o��o���? ��u5��E�k�}� �����)���M��� �1���U���ˏݏa� y��ӟ�I��m�� H���c�ǟ�������� !�3���W��{�'�M� ӯïկ�����/� ۿ��w�7ϛ����� 9�㿏ϵ���+���O� a�s���Eߩ�i�{��� ������9���]�� /��E��	���߭� ������Y��}�� �����q�������� 1�C�U�������K] ��i������? �u'��t $�S">/y� 3 �"y !��	
 �/�'/~�UD1:\4,����R_GRP� 1?;� 	 @� /�+{/@�/�/�/�/�/�.�	0  ?.:�!4/X?C?|?g5?�  �?�;�?�? �?�?�?O�?!O#O5O kOYO�O}O�O�O�O�O�O_	G!_3_��SCB 2@� �?_�_�_�_�_��_�_�_oUTORIAL A��/Zo�V_CON?FIG B�! �`/Ko�oog�OUTPUT yC��`���o 	-?Qcu��������a�)�\Regular� Option\�R713 : E�therNet/�IP Safety�4�F�X�j�|��� ����ď֏���o� �/�A�S�e�w����� ����џ��t��� � 2�D�V�h�z������� ¯ԯ���
��.�@� R�d�v���������п ����*�<�N�`� rτϖϨϺ������ ��&�8�J�\�n߀� �ߤ߶���������� "�4�F�X�j�|��� ������������0� B�T�f�x��������� �������,>P bt������ ��e��o�o4FX j|������ �/��0/B/T/f/x/ �/�/�/�/�/�/�/? /,?>?P?b?t?�?�? �?�?�?�?�?OO'? :OLO^OpO�O�O�O�O �O�O�O __#O6_H_ Z_l_~_�_�_�_�_�_ �_�_o_2oDoVoho zo�o�o�o�o�o�o�o 
-o@Rdv� �������� )<�N�`�r������� ��̏ޏ����%�8� J�\�n���������ȟ ڟ����"�3�F�X� j�|�������į֯����������>�P�:�)�{�)�\Regular� Option\�R713 : E�therNet/�IP Safety��ҿ�����,� >�P�b�t�'������� ��������(�:�L� ^�p߂�3��߸����� �� ��$�6�H�Z�l� ~�ߢ���������� � �2�D�V�h�z��� �����������
 .@Rdv���� ����*< N`r����� ��//&/8/J/\/ n/�/���/�/�/�/ �/?"?4?F?X?j?|? �?�/�?�?�?�?�?O O0OBOTOfOxO�O�? �O�O�O�O�O__,_�>_P_b_t_�_�^�$�TX_SCREE�N 1DR�;:��}��_�_ �_ oo$o6o�_�� �_vo�o�o�o�o�oGo Yo*<N`�o ��o������ y&��J�\�n����� ���-�ڏ����"� 4���X�Ϗ|������� ğ֟M���q��0�B� T�f�x�������ү �����,���P�b��t�������!�ο�$�UALRM_MS�G ?�Y��P ƿ�J ��C�6�g� Zϋ�~ϐϮϴ������	���-��SEV � �_�߲E�CFG F�U��Q  �E@��  A��   B)����P�к��h�� A!��Mh���ߒ�Mjs�q���MkFm~�� �Mm?s�߿o�MtP$� � .Mcgh� ��|2�H�jMc���N�sMdt�L6�ΖMfqF~k�GRP 2Gu�� 0�҃�	 ����@��ڂ�����:%����-���Y[�4�I_BBL_N�OTE Hu�T��l�B�P�A����DEF�PRO�%� �(%��IN.�L�% !�p�[���������� �� ��6!Z���FKEYDATA� 1I�Y  	�p �כF �d�����,�(9�D'OIN�T T>ACC�ANCE}��C	�PREV STE9P�DEXT��>}FINISM�/�� ORE INFO/ /]/o/V/�/ z/�/�/�/�/�/?#?�
?G?.?k?}? ���/frh/g�ui/white�home.png�~?�?�?�?�?O� } �5point�?�8OJO\OnO�OF/�FRH/FCGT�P/wzcancel'O�O�O�O�O	_zA�Jprev�O�C_U_g_y_�_E�Inex&O�_�_�_�_o��O�@finish��_Mo_oqo�o�o�]info<o�o�o�o G1CUgy� �,����	�� �?�Q�c�u�����(� ��Ϗ����)��� M�_�q�������6�˟ ݟ���%���I�[� m���������5��� ���)�;�B�_�q� ��������H�ݿ�� �%�7�ƿI�m�ϑ� �ϵ���V������!� 3�E���i�{ߍߟ߱� ��R�������/�A� S���w������� `�����+�=�O��� a�������������n� '9K]��� �����j� #5GYk���������;���0�0/B/�2/�k/}/�3,c?�/[8O?INT ER�/�/? IRECT�/?Ɨ ND�/1?`3CH�OICE]5?7? ?OUCHUPa?b? �?�?�?�?�?�?O�? /OOSOeOLO�OpO�O�O�O�O­frh/�gui/whitehome�o(_:_�L_^_p_�TUpoin�_�_�_�_�_�_~_i/direc�_ ,o>oPobotoo�`o��o�o�o�o�o�o
Qchoic_4FX�j|/touchup$����|��^arwrg�o <�N�`�r���{���� ̏ޏ�����&�8�J� \�n�����!���ȟڟ ������4�F�X�j� |������į֯��� ����B�T�f�x��� ��+���ҿ����� �O��P�b�tφϘϪ� ����������(߷� L�^�p߂ߔߦ߸�G� ���� ��$�6���Z� l�~����C����� ��� �2�D���h�z� ��������Q�����
 .@��dv�� ���_�* <N�r���� �[�//&/8/J/ \/��/�/�/�/�/�/ i/�/?"?4?F?X?/��f;��@����?�?�=�?�?�?�6,�OO�O<O#O`O rOYO�O}O�O�O�O�O �O_&__J_1_n_�_ g_�_�_�_�_�_�_�_ "o	oFoXo7�|o�o�o �o�o�o�/�o0 BTf�o���� ��s��,�>�P� b����������Ώ�� 򏁏�(�:�L�^�p� ��������ʟܟ�}� �$�6�H�Z�l�~�� ����Ưد����� � 2�D�V�h�z�	����� ¿Կ���
ϙ�.�@� R�d�vψ�ϬϾ��� ����ߕ�*�<�N�`� r߄ߖ�mo�������� ���8�J�\�n�� ���3���������� "���F�X�j�|����� /���������0 ��Tfx���= ���,�P bt����K� �//(/:/�^/p/ �/�/�/�/G/�/�/ ? ?$?6?H?�/l?~?�? �?�?�?U?�?�?O O 2ODO�?hOzO�O�O�Oh�O�O���K�������O_#]�OE_W_1V,Co�_;o �_�_�_�_�_o�_*o <o#o`oGo�o�o}o�o �o�o�o�o�o8 \nU�y���� ���"�4�F�UOj� |�������ď֏e��� ��0�B�T��x��� ������ҟa����� ,�>�P�b�񟆯���� ��ί�o���(�:� L�^���������ʿ ܿ�}��$�6�H�Z� l����Ϣϴ������� y�� �2�D�V�h�z� 	ߞ߰��������߇� �.�@�R�d�v��� �����������*� <�N�`�r�������� ��������8J \n��!��� ���4FXj |��/���� //�B/T/f/x/�/ �/+/�/�/�/�/?? ,?�/P?b?t?�?�?�? 9?�?�?�?OO(O�? LO^OpO�O�O�O�OGO �O�O __$_6_�OZ_ l_~_�_�_�_C_�_�_@�_o o2oDo�Fk�������oo�o�mko�o�o�f, ��o�@R9 v]������ ��*��N�`�G��� k�����̏ޏŏ�� &�8��\�n������� ���_ڟ����"�4� F�՟j�|�������į S������0�B�ѯ f�x���������ҿa� ����,�>�P�߿t� �ϘϪϼ���]���� �(�:�L�^��ςߔ� �߸�����k� ��$� 6�H�Z���~���� ������y�� �2�D� V�h������������ ��u�
.@Rd vM������� ��*<N`r� �����/� &/8/J/\/n/�//�/ �/�/�/�/�/?�/4? F?X?j?|?�??�?�? �?�?�?O�?0OBOTO fOxO�O�O+O�O�O�O �O__�O>_P_b_t_ �_�_'_�_�_�_�_o o(o�_Lo^opo�o�o �o5o�o�o�o $ �oHZl~���ڋ �{�� �������%�7��,#�h����s� �����͏
��� @�'�d�v�]������� П����۟���<�N� 5�r�Y������̯ޯ ���&�5J�\�n� ��������E�ڿ��� �"�4�ÿX�j�|ώ� �ϲ�A��������� 0�B���f�xߊߜ߮� ��O�������,�>� ��b�t������� ]�����(�:�L��� p�����������Y���  $6HZ��~ �����g�  2DV�z�� ������
//./ @/R/d/k�/�/�/�/ �/�/�/�/?*?<?N? `?r??�?�?�?�?�? �??O&O8OJO\OnO �OO�O�O�O�O�O�O �O"_4_F_X_j_|__ �_�_�_�_�_�_o�_ 0oBoTofoxo�oo�o �o�o�o�o�o,> Pbt��'�� �����:�L�^� p�����#���ʏ܏�� ��$��&��>����O�a� s�K�������,��؟ ����� �2��V�=� z���s�����ԯ�ͯ 
��.�@�'�d�K��� o��������ɿ�� �<�N�`�rτϖϥ� ����������&ߵ� J�\�n߀ߒߤ�3��� �������"��F�X� j�|����A����� ����0���T�f�x� ������=������� ,>��bt�� ��K��( :�^p���� �Y� //$/6/H/ �l/~/�/�/�/�/U/ �/�/? ?2?D?V?-� z?�?�?�?�?�?�/�? 
OO.O@OROdO�?�O �O�O�O�O�OqO__ *_<_N_`_�O�_�_�_ �_�_�_�__o&o8o Jo\ono�_�o�o�o�o �o�o{o"4FX j|����� ���0�B�T�f�x� �������ҏ���� ��,�>�P�b�t���� ����Ο������(��:�L�^�p�����k0����k0�����ѯ㭻����,�H���l�S����� ��ƿ������ �� D�V�=�z�aϞϰϗ� �ϻ������.��R� 9�v߈�g?�߾����� ����*�<�N�`�r� ���%��������� ���8�J�\�n����� !�����������" ��FXj|��/ �����B Tfx���=� ��//,/�P/b/ t/�/�/�/9/�/�/�/ ??(?:?�/^?p?�? �?�?�?G?�?�? OO $O6O�?ZOlO~O�O�O �O�O���O�O_ _2_ D_KOh_z_�_�_�_�_ �_c_�_
oo.o@oRo �_vo�o�o�o�o�o_o �o*<N`�o ������m� �&�8�J�\������ ����ȏڏ�{��"� 4�F�X�j��������� ğ֟�w���0�B� T�f�x��������ү ������,�>�P�b� t��������ο����@���@���/�A�S�+�uχ�a�,s߸�k��� �� ����6��Z�l� Sߐ�wߴ��߭����� � ��D�+�h�O�� �����������O� .�@�R�d�v������� ����������*< N`r���� ���&8J\ n��!���� �/�4/F/X/j/|/ �//�/�/�/�/�/? ?�/B?T?f?x?�?�? +?�?�?�?�?OO�? >OPObOtO�O�O�O9O �O�O�O__(_�OL_ ^_p_�_�_�_5_�_�_ �_ oo$o6o�Zolo ~o�o�o�o�_�o�o�o  2D�ohz� ���Q��
�� .�@��d�v������� ��Џ_����*�<� N�ݏr���������̟ [����&�8�J�\� 럀�������ȯگi� ���"�4�F�X��|� ������Ŀֿ�w�� �0�B�T�f����Ϝ� ��������s���,��>�P�b�t��$UI�_INUSER � �������  �u�y�_MENHI�ST 1J���  ( ��Є�'/SO�FTPART/G�ENLINK?c�urrent=m�enupage,/34,4��9��*��<�N���)�� �1133,1 OT�� ����������߃�� 3 _1,5��6�H�Z���(���48,2f�������������,18��LABEL���@Rd�o���5�N,8�n���c���631#��BTf��y-�edit��FIND_BOX`3�������� ��!/*/</N/`/r/�/ /�/�/�/�/�/ ?�/'?9?K?]?o?�? ?�?�?�?�?�?�?O �?5OGOYOkO}O�OO �O�O�O�O�O_�O1_ C_U_g_y_�_�_,_�_ �_�_�_	oo/?oQo couo�o�o�o�_�o�o �o)�oM_q ���6���� �%�7��[�m���� ����D�ُ����!� 3�W�i�{������� ßR������/�A� ,oJ�w���������ѯ ԟ����+�=�O�ޯ s���������Ϳ\�޿ ��'�9�K�]�쿁� �ϥϷ�����j���� #�5�G�Y���jߏߡ� ��������x���1� C�U�g�R� ����� ���������-�?�Q� c�u������������ ����);M_q ������ �%7I[m�  �����/��3/E/W/i/{/�/x���$UI_PANE�DATA 1L�����!�  	�}/�FRH/FCGT�P/FLEXUI�F.HTM?co�nnid=0 h�eight=10�0&_devic�e=TP&_li�nes=3� columns=4� �fon� 4&_p�age=doub�� 1�/v�)prsim=?f?  }i?��?�?�?�?�?�? ) �?O�?1OOUOgONO��OrO�O�OL110q7�O�OL195�O�_K2
SYSVA�RS.SV  A�ME.TP_}�ߐ� _P ���nw4fr�h/cgtp/f�lex� .stm�?_width=�� �/02??*62I_�Hual�_om[itree�Q	oAo Soeowo�_�o�o�o�o �o�o�o+Oa H�l����RX� � _P  ா!{? �2� D�V�h�z����q? ԏ���
����@�R� 9�v�]�������П�� ��۟�*��N�5�r����u���#����ү �����m�>���b� t���������#��� ٿ���:�L�3�p�W� ��{ϸ��ϱ������ $ߗ���Z�l�~ߐߢ� �����K���� �2� D�V�h��ߌ�s��� ������
���.�@�'� d�K���������1�C� ��*<N��r ��ߨ���� i&J\C�g ������/� 4//X/������/�/ �/�/�/�/M/?�B? T?f?x?�?�??�?�? �?�?�?O,OOPO7O tO[O�O�O�O�O�O�O _w/�/:_L_^_p_�_ �_�O�_+?�_�_ oo $o6oHo�_loSo�owo �o�o�o�o�o  D+hza�_#Z������*�<�)�a��UP������� ÏՏ�N���/�� (�e�L���p������� �ʟ�� �=��X'S�![�$UI_PO�STYPE  �'U� 	� �qI��Zo�Q�UICKMEN ; ~� �����_RESTOREw 1M'U����*de�fault�[�DOUBLE��PRIM�m�menupage?,153,1J�}�P������V�^�3i� �����R�*�N�`� rτϖ�)�0��Ϲ�+� ����*�<�N���r� �ߖߨߺ�]������ �&���3�E�W��ߒ� �������}����"� 4�F�X���|������� ��o�������g�0B Tfx���� ��,>P�� o������ //�:/L/^/p/�/�%/�/�/�/�/�/��S�CRE��?í�u1sc��u2/43/44/45*/46/47/48/13wTATz�� ң<'Ug�USER0?�(4ks13�43�44��45�46�47�48��1o�NDO_CFOG N~���o��PDr1�9��None���0_INFO 1O'U5V@Р0%�/qO �X_O�O�O�O�O�O�O _�O0__T_f_I_�_��__�_��CAOFF?SET R~�ZA�_�#��/o#o5o Gotoko}o�o�o�o�_ �o�o:1Cp gy��kӯ�}���
���XUFRA�M3��$F@AR�TOL_ABRT8C�>C[�ENBd�U�?GRP 1S�ϡCz  A��� ��A��ʏ܏� ��$�6�W���U��As�?MSK  ��VAi���W�N@�%NI��%FIND_�BOX&���VARS_CONFI@�T�[ FP�#�n֘CMR��2Z�['h�� 	@����P1: SC130EF2 *S��W��$��h������5� A?�F�@�F�p:��̞ ������(֯���:��=���4�A��")�z��" B��͕��!��!� ���޿����&�� J�5�Gπ�׿a϶ϡ�����ϟ��"�ڔISIONTMOUc����E�9�B�[�x��䯁 FR:�\;�\$@A\'� �� MCz��LOG��   7UD1z�EX�ߗ!�' B@ ���ҿѧ����4�# � n6  ����&���j��`F�С?  =��͂�$������TRAI�N��J���  d���p��o�Z��\�](����
����� '�9�K���o����������������#��9�_��REe�]��@�ڔ/LEXEb�^�@�1-=@ОMPHA%St0+EC��ۓ�RTD_FILT�ER 2_�[ ��eȢ��+ =Oas���j� ����/"/4/F/�X/j/ؖSHIFT�a�1`�[
 <��%���/�4�/�/? �/�/8??!?n?E?W? }?�?�?�?�?�?�?"O��?	LIVE/�SNA��%vs�fliv�4O��;� �PU��WBmenumOrOO�O�O��B�%b�a�)t�%M�Ob�bt�E��$�WAITDINE#NDF�p�CTO��g��aWD�w_S�_^YTI]M�����\GH_ �]j_�[�_�Z�_�Z�_\XRELE���@T�Aߑ�,AS_AC�TJ@�h��]W_�� �c��:�AN_S�LOc�+��bRD�IS�����$XS�c�d��~�/���EpV�Rc�et�$Z�ABC��fQ �,�2*�ZIPb�gQ���$��6��zMPCF_Gw 1h�� 0�����N��si_����� ���֏��<x�ۏ��ŏ:�� ����Y�?�)���M�o� ş����
��ſ��%� �1�G�U���pW�e��j��s�pYLINuD�k_� �M�,(  *����`ݯ��>�%� � t�����گ��*�߿ƿ ؿ�X�9�K�]Ϡ��� �ϷϞ�����0�ߘ#��{��2l_��a �t�n�~�gs��@����ϙ^���ϗ���A���SPHER/E 2m���u�Q� ��J��n������� ��o�����M�4�q� X������ ����b� ��I��m�6�pZZ�f Ǖf