��   �A��*SYST�EM*��V9.1�060 11/�14/2017 A 	  ����HAPTIC�_T   8 �$ENABLE�  $BBLNOTEENB=�MAX_ALAR�MSLIO=��4&ALM- � $ERRCsOD<' STY;�kIO- X ��
$IOTYP�<$INDEX��TRG�RSR;V1�VAL=��2�3=�HPC�FG- $ �6$DEBUG�=COMP_SW���$$CLAS�S  ����C��f��f8VE�RSION@�  �����* / af���l�
�r_D�F� 2C��(   �� #�5��V�C�D�2 \������/./@/R/d/v/ �/�/�/�/�/�/��MF�   `�<	"T�9G��C�G��;284`8 @9x?�?�?�?�?�?�?H�?�d 2?6�
  +O=OOOaOsO�O�O�O@�O�O�O�O_�+Uu ">
	/K_]S�3U���_�_�_�_�%P_�MOT_	C ��R