��   9�A��*SYST�EM*��V9.1�060 11/�14/2017 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG4��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST��wNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !�� FT� @�� LOG_8	,C�MO>$DNL�D_FILTER��SUBDIRCAPCΌ �8 .� 4� H{A�DDRTYP�H NGTH���4�z +LSq� D $ROB�OTIG �PEEyR�� MASK��MRU~OMGD�EV�gPINF�O�  $�$$TI ��RCM+T� A$( /�QS�IZ�!S� TA�TUS_%$MA�ILSERV �$PLAN� <�$LIN<$C�LU��<$TOޥP$CC�&FR\�&YJEC|!Z%�ENB � ALkAR:!B�TP,��#,V8 S��$�VAR�)M�ONx�&���&APPL�&�PA� �%��'PO�R�Y#_�!�"AL�ERT�&i2URL� }Z3ATT�AC��0ERR_oTHROU3US�9H!�8� CH- c%�4wMAX?WS_|1w��1MOD���1I�  �1o (��1PWD  � L�A��0�ND�1T{RYFDELA-Cx�0G'AERSI���1Q'ROBICLK�_HM 0Q'� XML|+ 3SGFRMU3�T� !OUU3 G_�-COP1�F33ĿAQ'C[2�%�B_A�U�� 9 R�!U{PDb&PCOU{!��CFO 2 �
$V*W�@c%AsCC_HYQSNA�_UMMY1oW2?_4�RDM* �$DIS�S=M	 l5��o!�"%Q7�IZP�%H� �VR�0�UP� �_DLVSPAR���QN,#
3 ��_�R!_WI�CT?Z_INDE�3^`gOFF� ~URmi�D�)c�  � t Z!`MO�N��cD��bHOUU#E%A�f�a�f�a��fLOCA� #{$NS0H_HE�K��@I�/ 3 �$ARPH&�_7IPF�W_* O2�F``QFAsD90�VHO_� 5Rr;EL� P��r�90WORA5XQE� LV�[:R2�ICE��p����$cs  �����q��
��
��p�PS�A�w�  ���$X'0 
�
���F������F�?��$.� 2'��r����rw�X��� '���!��q�����$� _F�LTR  	�2�� ���������ы$'�2ы7rS�H`D 1'�" P��o�<�^��� ������㟦��ʟ� �<�a�$���H���l� ͯ��񯴯Ư'��K� �o�2���V�h�ɿ�� ���Կ5���.�k� ZϏ�Rϳ�v��Ϛ��� ���1���U��y�<� ��`��߄ߖ��ߺ�� ��?��c�&�8��\� �����������;��*�_�"���Շz _L�UA1�x!1E.��0��F���1��>F�255.��&H��D���2����@: ����13;���� as��14 ���*���15+���Qcu�16��� �����I��Q��������h�X�|�� 'Q� {�K.<�/�/ �/�/ ?2?D??h?z?C�PY?�?�?�?�?�? OO(O�?LO^OpOK.�AOB�G��O�L
�ZDT Status0O�O__/_D��}iRConn�ect: irc�QT//alert �Nz_�_�_�_CW�O�_@�_oo&o8oJ�4�PT2=���=oso�o �o�o�o�o�o�o�'9KB�$$c9�62b37a-1�ac0-eb2a�-f1c7-8c�6eb5418bb9  (�_��O ����F�!-��(�")��J�� 0.��C� }�,$�v� -���d�����ŏ��ҏ �����C�U�<�y� `�������ӟ����ޟ�K�(���� D�M_�!����S�MTP_CTRLg 	��u�%� ���D�p���J�ٯ�į���LP�NU��!
�@��O�G�!����\n�Ԉ#"�US?TOM @�i��r��  r�$T�CPIP:�@���H�%��TEL������!�h�H!T�Vb�D�rj3/_tpd� ��?�?!KCL���?�q��!CRT�x�fϿϣ"G�!OCONS���-�ib_smon����