��   ��A��*SYST�EM*��V9.1�060 11/�14/2017 A   ������DMR_S�HFERR_T �  $O�FFSET  � 	4/GR�P:� $�MA��R_DON�E  $OT�_MINUSJ � 	sPLzdC�OUNJ$REF,j�PO{���I$BCKLSH�_SIG�EA�CHMSTj�SsPC�
�MOVn �~ADAPT_I�NERJ FR�ICCOL_Pz,MGRAV��� HISID�SPk�HIFT�_7 O �N\m�MCH� S��ARM_PARA�O dcANG�o y2�CLD�E7�CALIB�Dn$GEA�R�2� RING,��<$]_d��REL3� 1  	4�CLo�: � �A�X{  $PS_��TI���TI�ME �J� _gCMD��"FB��VA �&CL_OV��� FRMZ�$DmEDX�$NA� �%�CURL��W���TC�K�%�FMSV��REM_LIF	��'83:c$,�-9_09:_��=��%3d6W� �"�P�CCOM��FB� M�0�MAL_F�ECI�P:!no"DTYkR_|"8�5:#�1END�4�y�o1 P sPL� W ���STA:#TRQ_�M��� KNYFSD� eHYcJ� XGIpJuI~JI�D4�$��ASS> �����A�����@VE�RSI� �G�  ���$�S 1�H ���� 	 ���.__R_=Vw�D |�� Ɇ������ �" ��Y_C_�_ �_�_�_���@�R�_�C�ol�� (�  6�HyP�� i�J��> obo�_'l�o�o�o�o��`��!� �M�� �@�oUiO @Btp
u@�o_oH3l��d_�����=L�����?����@� �4�F�X�j�|��������ď֏���M ��E%�3��S��D  2���������̟ޟ ���&���<s�P� b�t���������ί�@������@D�(] J�Yn�Y���}����� ���׿���4��X��C�hώ��$4 1�\�y�M���KZ:�L�q�)F�5UV��oO�K�m�E����G��ED��G�9}�y<G���?a�m�B���k���ZH���D���nӸ�e�+¨�CC��d��ҖhH�5E"��:��= ?�B�m�oAɒ��ߒ�m�*�������-����Me�y���u�����3����My�F�M{@�*��A��� �G�M�x56�OY	A�������?��>d©��B���*�OYA�������?���©��B���b�:=�O��U����6�ҩ�=������2  ��%T?OTESCA�e&��������W6�I��=AA�6����P?�gv¦埬B���9�V�B�AA�9�����?���¦���B���9���:2�Z��q;����߻�_�;����a���1�C���R��A@ԣ����^?��\¦?g�B���n������ժ?��Z�¦��B���@9�������0L�����@\ O>�oΠ�������F��R���A<�����?��£���B��<.���A<����?�~�¤�B������p���>i��:�ާ����~�a��F�\��2��@W*������?���«��B�x\�2���@WV������?��O«S~��>  �%�����<3t �mg�	��>�P!/t�B/6���f��%b���4�?{��¤���C!����f��%x������?|\¤�ȔC!m� � ��Z������<s >N������/�/4/F��-�R#J�� ��M��&�?{�o�¦^�j ��n/J�� ���� ?{�����C!p9����������x�rA ������_a�P�&DEMaO�/�?5�:�T6��EH�����=~�{�D���B�sR��E��	N�����zǨ��TB�z�V>������ U;��sJ%�z�(�?hO�B�
|�6��-Z������²)����¨=BC�8���A�����ؾ�6§��gC�L�/  ��^�+?��,��!V�@ۮGo���>O��"VIZPIXoO��B�h16ҽ�o��������>��K¥��mC�����o����@�U����Y¦I�Cէ9��I��3�	��E��̼`x�@]��?���a�Q�_��_�$B\6RT�������z����¥��C���n_p����Y�ݳ����¦ lC���9�<7��������
����@��?��2�^�_�_�o�%B[p�b6������{�^������6�¥��C�����c��������r8��y����4C��V���ي���j���x�A��A�R�~~o�oa4_�F�Qd9J������u�����¦��C���.o9[��O�k���m�� �O§%Cy�H9��Z����^��F>���A��o���z�>P!�t�wn��6Ҿ��F!���N�����H¯��BZ��������FN����(C��\��¯�qB[�b�O=֔�߾JQD;��� ����ޏ�?�C���:���5����zU�e��¨�]N�U�V����T�9h��¨�C����O  �]3I߿��S;�$'�p��g�/ ��  �%MA!I�/����6�u v% Viޟt'����0�~� �h_��mVg̟����� ��ί��J��-���� `�N���r������� 4�F������J�8�n� Ŀֿ�������X��π���4ߊ�[�m�����$PLCL_GR�P 1%��� D&�?�  ����*���&�	� ��-��Q�<�N��r� ������