��   ,��A��*SYST�EM*��V9.1�060 11/�14/2017 A   ����DCSS_I�OC_T   �P $OPER�ATION  $L_TYPB7IDXBR1H[ �S2]2R4�$�$CLASS  �������Pz��P� VERS?��  ����$' 2 ��P @� ������
H�� ����� ����"� "I[m��� ����/!/3/E/ W/i/{/�/�/�/�/�/ �/�/??/?A?S?e? w?�?�?�?�?�?�?�? OO+O=OOOaOsO�O �O�O�O�O�O�O__ '_9_K_]_o_�_�_�_ �_�_�_�_�_o#o5o GoYoko}o�o�o�o�o �o�o�o1CU gy��������_C_CCL ?���  	�All para�m��
Base��Pos./�Speed ch�eck(�Safe� I/O con/nect�}R��`� �2�D�V�SIi��@{�exter�nal_esto�p����fence ���'�9�K�b�o��� ������ɟ۟���� #�:�G�Y�k������� ��ʯׯ�����1� C�Z�g�y��������� ӿ���	��2�?�Q� c�zχϙϫ������� ��
��)�;�R�_�q� �ߚߧ߹�������� �*�7�I�[�r��� �������O�{��auto_di�sabled��in ���C�U�~�y� ������������	 -VQcu�� �����.) ;Mvq���� ��///%/N/I/ [/m/�/�/�/�/�/�/ �/�/&?!?3?E?n?i? {?�?�?�?�?�?�?�? OOFOAOSOeO�O�O��O�O�O�O�O�� �N�  ���	_��;_ M___q_�_�_�_�_�_ �_�_oo%o7oIo[o moo�o�o�o�o�o�o �o!3EWi{ ����������SIh���#��f� x���������ҏ��� ��,�>�P�b�t��� ������Ο����� (�:�L�^�p������� ��ʯܯ� ��$�6� H�Z�l�~�������ƿ ؿ���� �2�D�V� h�zόϞϰ������� ��
��.�@�R�d�v� �ߚ߬߾����������*�5�P%_�SOFDI10�y�2�y�3��y�4��y�5$��y�6��y�7��y�8�G�3�E�W�n�{� �������������� /FSew�� �����+ =Ofs���� ���//'/>/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?^?k? }?�?�?�?�?�?�?�?@OO6OCON�`�Od�v�O~�C��C��C ��C��C��C��C &�A�Q_c_�_�_�_�_ �_�_�_�_oo)o;o do_oqo�o�o�o�o�o �o�o<7I[ ������� ��!�3�\�W�i�{� ������Ï����� 4�/�A�S�|�w����� ğ��џ����+��T�O�a�lO_�Sc��v�VOFFn�F�ENCE��EX�EMGկ���N�TED�OP���AUTO��T�O[��O�M�CC|��CSBP���
POSSP�D_ENB�C�ONF_OK��F�_IPAR_CR(�����Ov�_๯Bձ_Я;���'��DIS��C_D���_`���y� 