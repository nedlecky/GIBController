��  Ij�A��*SYST�EM*��V9.1�060 11/�14/2017 A   ����SBR_T �  | 	$S�VMTR_ID � $ROBO�T9$GRP�_NUM<AXIaSQ6K 6NFF�3 _PARAM�F	$�  �,$MD SPD�_LIT4&2�*  � ���4�$$C�LASS  ����������� VERSION��  ����$'  1 ~� T����M-10iA�_Enh_Wri�st���  �aiS8/400�0 40A��
�H1 DSP1-�S1��	P01�.0e,  �	�  ��
PCR ��} �C������0��{  ����r9�  3!M�����  �H�  �����
/�m���  X���< �mm��  ����R �2.h��>�����7(��h�����&���
= �b ���� �6����������g 2 �g���"2����.����B�� � d ���c �8 �:?����'b:
�@E/�/�/�/�/���?��f?C?U?g?���2D+�
 ������g^�2�&�
 �<�"���a?p?�?���0BT2b^2fx��P����������W 5�/7�/7��@��?� 3!���=��y��p��c5\�+�Z, r ���4 /8$��?����d O\/��r(�~/�/rD�/r_ �_�_�_?�_'?�_o�o&o 4�����<]����W���1��1=��>���� ?G2(oso���t�?2�22/5A�2O3^3O0N��  8@��������{���bD�<��9"�R8� l� �� �&��3�Pp�9S9� � ���}3�(YR`^��N p� �?�Y�+:@= � ��� �<8$�zosC � mjS������� ��Or(��c9	`t �# (��� ���LTqTYa��-�?�Q�c��_�� �_����Ϗ�����)���@�o0�biS0.5/)6�kZ4^4�o0M���� ��_�Kn���Hw�HbD����&s(p �8 �����v�|� x����5@#�5���� ��� +8$�pi�n�rB��S�DP���utC�P�%}����s�p2�:���!�TY��~���
	m� ���r�;���_�q����������˿ݿ�:�\F�0l�Ro��Z5^�A��������~��, �p�~�<<؟� -��{� ��������� � �r-��r� �Sp�����e��r(M����ʯܯ�߷� ��$���H���#�5�G�`Y�k�}������*0"�4+�6^7"�J�4G@Ah�d�R��ax�3��t��a�8	�k�����0�;L� ����������� 7 ���� p8$���5b� gZ�S������ׇ�y����s�tf�xАTY �r>���)���c u��߫������"4FX �����ZP��on0g�	�V�����// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?2<�2?V?h?z?�?�?�? �?�?�?�?
OC�~ (O����O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_�_ @?oo,o>oPoboto �o�o�o�oOJO<O `OrO:L^p�� ����� ��$� 6�H�Z�l�~����_�� Ə؏���� �2�D� V�h�z��o���� 0��
��.�@�R�d� v���������Я��� ��*�<�N���r��� ������̿޿��� &�8ϴ���P�ʟܟ� �����������"�4� F�X�j�|ߎߠ߲��� �������h�0�B�T� f�x���������� @�r�d�-��Ϛ�b�t� �������������� (:L^p�� ����� $ 6HZl~���� ��4�F�X� /2/D/ V/h/z/�/�/�/�/�/ �/�/
??.?@?R?d? v?��?�?�?�?�?�? OO*O<ONO`O�� xO�//�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o �?Xojo|o�o�o�o�o �o�o�ohO�O�OU �O�O������ ���,�>�P�b�t� ��������Ώ��<o� �(�:�L�^�p����� ����ʟ&��\n �H�Z�l�~������� Ưد���� �2�D� V�h�z�������¿Կ ���
��.�@�R�d� vψ�������,�>� ��*�<�N�`�r߄� �ߨߺ��������� &�8�J�\︿���� �����������"�4� ���ϴ�}����ϲ��� ������0BT fx������ �d�>Pbt �������N� /
/������p/�/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�? �?"�?�?O O2ODO VOhOzO�O�O�O,// �OB/T/f/._@_R_d_ v_�_�_�_�_�_�_�_ oo*o<oNo`oro�o �?�o�o�o�o�o &8J\�O�O�O�  __����"�4� F�X�j�|�������ď ֏�����0��oB� f�x���������ҟ� ����v?�2��� �������ί��� �(�:�L�^�p����� ����ʿܿ�J��$� 6�H�Z�l�~ϐϢϴ� ����T�F���j�|��� V�h�zߌߞ߰����� ����
��.�@�R�d� v����������� ��*�<�N�`�r��� ������(�:� &8J\n��� �����"4 FX��j���� ���//0/B/�� g/Z/�������/�/�/ �/??,?>?P?b?t? �?�?�?�?�?�?�?O Or:OLO^OpO�O�O �O�O�O�O�O _|/n/ _�/�/�/~_�_�_�_ �_�_�_�_o o2oDo Vohozo�o�o�o�o�o 0O�o
.@Rd v���_:_,_� P_b_*�<�N�`�r��� ������̏ޏ���� &�8�J�\�n����o�� ��ȟڟ����"�4� F�X�j��������  ������0�B�T� f�x���������ҿ� ����,�>Ϛ�b�t� �ϘϪϼ�������� �(ߤ���@ߺ�̯ޯ �߸������� ��$� 6�H�Z�l�~���� ��������X� �2�D� V�h�z����������� 0�b�T�xߊ�Rd v������� *<N`r� ������// &/8/J/\/n/�/�/�� �/�/$6H?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fO��O�O�O�O�O�O �O__,_>_P_�/�/ h_�/�/?�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ �OHZl~��� ����X_�_|_E� �_�_z�������ԏ ���
��.�@�R�d� v���������П,� ��*�<�N�`�r��� �������߯үL�^� p�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώ�ꟲ��� ��������0�B�T� f�x���毐�
��.� ����,�>�P�b�t� ������������ �(�:�L���p����� ���������� $ �߲ߤ�m���ߢ� ���� 2D Vhz����� ��T�
/./@/R/d/ v/�/�/�/�/�/�/> ?�/t��`?r?�? �?�?�?�?�?�?OO &O8OJO\OnO�O�O�O �O/�O�O�O_"_4_ F_X_j_|_�_�_?? �_2?D?V?o0oBoTo foxo�o�o�o�o�o�o �o,>Pbt �O������� �(�:�L��_�_�_�� �_oʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟���� �|2� V�h�z�������¯ԯ ���
�f�/�"����� ����������п��� ��*�<�N�`�rτ� �ϨϺ�����:��� &�8�J�\�n߀ߒߤ� ����D�6���Z�l�~� F�X�j�|������ ��������0�B�T� f�x������������� ��,>Pbt ����߽�*�� (:L^p�� ����� //$/ 6/H/��Z/~/�/�/�/ �/�/�/�/? ?2?� W?J?����?�?�? �?�?
OO.O@OROdO vO�O�O�O�O�O�O�O _b/*_<_N_`_r_�_ �_�_�_�_�_�_l?^? o�?�?�?no�o�o�o �o�o�o�o�o"4 FXj|����  _����0�B�T� f�x������_*oo� @oRo�,�>�P�b�t� ��������Ο���� �(�:�L�^�p���� ����ʯܯ� ��$� 6�H�Z����r���� �ؿ���� �2�D� V�h�zόϞϰ����� ����
��.ߊ�R�d� v߈ߚ߬߾������� ���0謹��ο ������������ &�8�J�\�n������� ��������H�"4 FXj|����  �R�D�h�z�BT fx������ �//,/>/P/b/t/ �/�/���/�/�/�/? ?(?:?L?^?p?�?� �?�?&8 OO$O 6OHOZOlO~O�O�O�O �O�O�O�O_ _2_D_ V_�/z_�_�_�_�_�_ �_�_
oo.o@o�?�? Xo�?�?�?�o�o�o�o *<N`r� �������� p_8�J�\�n������� ��ȏڏ�Hozolo5� �o�oj�|�������ğ ֟�����0�B�T� f�x����������ү ����,�>�P�b�t� �������Ͽ¿<�N� `�(�:�L�^�pςϔ� �ϸ������� ��$� 6�H�Z�l�~�گ�ߴ� ��������� �2�D� V�h��ֿ������ ����
��.�@�R�d� v��������������� *<��`r� ������ p���]����� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/D�/?0?B?T? f?x?�?�?�?�?�?. �?�?dv�PObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_?�_�_�_ oo$o 6oHoZolo~o�oO�? �o"O4OFO 2D Vhz����� ��
��.�@�R�d� �_��������Џ�� ��*�<��o�o�o�� �o�o��̟ޟ��� &�8�J�\�n������� ��ȯگ����l�"� F�X�j�|�������Ŀ ֿ���V��ό��� ��xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼���*���� �(�:�L�^�p��� ���4�&���J�\�n� 6�H�Z�l�~������� �������� 2D Vhz��߰�� ��
.@Rd ���������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?�J?n?�?�?�? �?�?�?�?�?O"O~ GO:O����O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_�_ �_R?o,o>oPoboto �o�o�o�o�o�o\ONO �orO�O�O^p�� ����� ��$� 6�H�Z�l�~������� o؏���� �2�D� V�h�z����o՟ 0B
��.�@�R�d� v���������Я��� ��*�<�N�`���r� ������̿޿��� &�8�JϦ�o�b�ܟ�  ����������"�4� F�X�j�|ߎߠ߲��� ��������z�B�T� f�x���������� �����v� ��ϬϾ� �������������� (:L^p�� ����8� $ 6HZl~��� �B�4��X�j�2/D/ V/h/z/�/�/�/�/�/ �/�/
??.?@?R?d? v?�?��?�?�?�?�? OO*O<ONO`OrO� �O�O//(/�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o Fo�?jo|o�o�o�o�o �o�o�o0�O�O H�O�O�O���� ���,�>�P�b�t� ��������Ώ���� `o(�:�L�^�p����� ����ʟܟ8j\%� ��Z�l�~������� Ưد���� �2�D� V�h�z��������¿ ���
��.�@�R�d� vψϚ����ϲ�,�>� P��*�<�N�`�r߄� �ߨߺ��������� &�8�J�\�n�ʿ��� �����������"�4� F�X�����p������ ������0BT fx������ �,��Pbt �������/ `�����M/�����/�/ �/�/�/�/�/ ??$? 6?H?Z?l?~?�?�?�? �?�?4�?O O2ODO VOhOzO�O�O�O�O/ �O�OT/f/x/@_R_d_ v_�_�_�_�_�_�_�_ oo*o<oNo`oro�o �o�?�o�o�o�o &8J\n��O�O �_$_6_��"�4� F�X�j�|�������ď ֏�����0�B�T� �ox���������ҟ� ����,����u� ������ί��� �(�:�L�^�p����� ����ʿܿ� �\�� 6�H�Z�l�~ϐϢϴ� ������F���|��� ��h�zߌߞ߰����� ����
��.�@�R�d� v���������� ��*�<�N�`�r��� ����$����:�L�^� &8J\n��� �����"4 FXj|���� ���//0/B/T/ �������/��
�/�/ �/??,?>?P?b?t? �?�?�?�?�?�?�?O O(O�:O^OpO�O�O �O�O�O�O�O __n/ 7_*_�/�/�/�_�_�_ �_�_�_�_o o2oDo Vohozo�o�o�o�o�o �oBO
.@Rd v�����L_>_ �b_t_�_N�`�r��� ������̏ޏ���� &�8�J�\�n�������  ȟڟ����"�4� F�X�j�|��
��ů  �2�����0�B�T� f�x���������ҿ� ����,�>�PϬ�b� �ϘϪϼ�������� �(�:ߖ�_�R�̯ޯ �������� ��$� 6�H�Z�l�~���� ���������j�2�D� V�h�z����������� ����t�f��ߜ߮� v������� *<N`r� ����(��// &/8/J/\/n/�/�/�/  2$�/HZ"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO��O�O�O�O�O �O__,_>_P_b_�%��$SBR2 1��%�P T0 �  @�/�' �_�_�_�_oo &o8oJo\ono�o�o�o �o�Q�o�_�o& 8J\n���� ���o��o"�4�F� X�j�|�������ď֏ �����0��T�f� x���������ҟ��� ��,�>�!�b�E��� ������ί���� (�:�L�^�p�S���w� ��ʿܿ� ��$�6πH�Z�l�~ϐϢυ�~ i_��������'�9� K�]�o߁ߓߥ߷��� �ظ���
��.�@�R� d�v��������� ������*�<�N�`�r� �������������� &
��\n�� ������" 4FX<f��� ����//0/B/ T/f/x/�/n�/�/�/ �/�/??,?>?P?b? t?�?�?�?�?�/�?�? OO(O:OLO^OpO�O �O�O�O�O�O�O�?_ $_6_H_Z_l_~_�_�_ �_�_�_�_�_o o_ DoVohozo�o�o�o�o �o�o�o
.@R 6ov������ ���*�<�N�`�r� ��h����̏ޏ��� �&�8�J�\�n����� ������ڟ����"� 4�F�X�j�|������� į֯��̟��0�B� T�f�x���������ҿ ������>�P�b� tφϘϪϼ������� ��(�:��^�p߂� �ߦ߸������� �� $�6�H�Z�l�Pߐ�� ����������� �2� D�V�h�z��������� ������
.@R dv������� �*<N`r �������/ �&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?/X?j?|?�?�?�? �?�?�?�?OO0OBO TO8?J?�O�O�O�O�O �O�O__,_>_P_b_ t_�_jO|O�_�_�_�_ oo(o:oLo^opo�o �o�o�o�_�o�o  $6HZl~�� �����o� �2� D�V�h�z������� ԏ���
�� �@�R� d�v���������П� ����*�<�N�2�r� ��������̯ޯ�� �&�8�J�\�n���d� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B� T�f�xߊߜ߮����� ������,�>�P�b� t����������� �����:�L�^�p��� ������������  $6�,�l~�� ����� 2 DVhLv��� ���
//./@/R/ d/v/�/�/~�/�/�/ �/??*?<?N?`?r? �?�?�?�?�?�/�?O O&O8OJO\OnO�O�O �O�O�O�O�O�O�?"_ 4_F_X_j_|_�_�_�_ �_�_�_�_oo0o_ Tofoxo�o�o�o�o�o �o�o,>Pb Fo������� ��(�:�L�^�p��� ��x��ʏ܏� �� $�6�H�Z�l�~����� ���������� �2� D�V�h�z�������¯ ԯ�ʟܟ�.�@�R� d�v���������п� ������&�N�`�r� �ϖϨϺ�������� �&�8�J�.�n߀ߒ� �߶����������"� 4�F�X�j�|�`ߠ�� ����������0�B� T�f�x����������� ����,>Pb t�������� (:L^p� ������ // �6/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?(/h?z?�?�?�?�? �?�?�?
OO.O@ORO dOH?Z?�O�O�O�O�O �O__*_<_N_`_r_ �_�_zO�O�_�_�_o o&o8oJo\ono�o�o �o�o�o�_�o�o" 4FXj|��� �����o�0�B� T�f�x���������ҏ �����,��P�b� t���������Ο��� ��(�:�L�^�B��� ������ʯܯ� �� $�6�H�Z�l�~���t� ��ƿؿ���� �2� D�V�h�zόϞϰ��� ������
��.�@�R� d�v߈ߚ߬߾����� �����*�<�N�`�r� ������������ ���
�J�\�n����� ������������" 4F*�<�|��� ����0B Tfx\���� ��//,/>/P/b/ t/�/�/�/��/�/�/ ??(?:?L?^?p?�? �?�?�?�?�?�/ OO $O6OHOZOlO~O�O�O �O�O�O�O�O_�?2_ D_V_h_z_�_�_�_�_ �_�_�_
oo.o@o$_ dovo�o�o�o�o�o�o �o*<N`r Vo������� �&�8�J�\�n����� ���ȏڏ����"� 4�F�X�j�|������� ğ��������0�B� T�f�x���������ү ���ڟ�,�>�P�b� t���������ο�� ��(��6�^�pς� �Ϧϸ������� �� $�6�H�Z�>�~ߐߢ� ����������� �2� D�V�h�z��p߰��� ������
��.�@�R� d�v������������� ��*<N`r ��������� &8J\n�� ������/"/ F/X/j/|/�/�/�/ �/�/�/�/??0?B? T?8/x?�?�?�?�?�? �?�?OO,O>OPObO tOX?j?�O�O�O�O�O __(_:_L_^_p_�_ �_�_�O�O�_�_ oo $o6oHoZolo~o�o�o �o�o�o�_�o 2 DVhz���� ���
��o.�@�R� d�v���������Џ� ���*�<�N�