��   X�A��*SYST�EM*��V9.1�060 11/�14/2017 A   ����CIPS_C�FG_T   �0 $INTE�RFACE  �$DUMMY1�B2B3B&SE�T/ @ $�MODA8 _S�IZ}OUT�DATE_FIX~�CSI_VRC �  4��$$CLASS ? �������O��O� VERS�ION�  ���$'1 �O� �m �r �
���  )) ,@