��   ��A��*SYST�EM*��V9.1�060 11/�14/2017 A   ����PMC_CF�G_T   �� $'NUM_�MSK  $�EXE_TYPE�CMEM_OPT�PN_CNFCI�F_CY:gSC�N_TIME �E RESET_PȂDo LJ �HECK_DSBLC �$DRA> AR�GINCSTOR�J�4&DEV�. d 	7O�C'HAR�AD�D�SIZORA�CBSLO[OD�KIOKOCCP�YC&l /  L ��h99�IDXC�L.o � 
�EQP�LHRAT�TRKBUF| ���UN_STATU�S�CU��MA�X(I��SNP�_PA�  �� � ANNE��� OW CTIO�N_�PU� �  $BAU}D�NOISYm�N�T1�#2�#3n�$_PR�T4P�' DATA�CQ�UEUE� PTH�[$MM_��%&!R�ETRIESCAUTO!R[���BG � �ISP_INFd�' C�LIMI� B5AD_H C3H��#d6�# d6�#d6�#W1� �#�4��#�4�#�4�"� �$�$CLASS  �����1��z���0VERSg ��8  7���iFG0 �5���
@+AT�2������d���3CC�  2G'@d $)DxO��uO �O�O�O�O�O�O__ :_)_^_M_�_q_�_�_ �_�_�_�_oo6o%o ZoIo~omo�o�o�o�o �o�o�o2!VE zi������ 
��.��R�A�v�e� ���������я��� *��N�=�r�a����� ����ޟ͟��&�� J�9�n�]��������� گɯ���"��F�5� j�Y���}�����ֿſ �����B�1�f�U� ��yϮϝ��������� �	�>�-�b�Q߆�u� �ߙ��߽������� :�)�^�M��q��� ���������6�%� Z�I�~�m��������� ������2!VE zi������ 
�.RAve ������/��*//N/=/R,CIFw 2aKP ^/ X/�/�/�/�/�/?? (?:?c?^?p?�?�?�? �?�?�?�? OO;O6O HOZO�O~O�O�O�O�O �O�O__ _2_[_V_ h_z_�_�_�_�_�_�_ �_
o3o.o@oRo{ovo �o�o�o�o�o�o *SN`r�� ������+�&� 8�J�s�n��������� ȏڏ����"�K�F� X�j���������۟֟��v/TYPE 2��+ (�R�d���L���"��h����������̠�����~#S�NP_PARAM' �+����  'C�q��@R���ݢQ�����UD�R�����