��   D�A��*SYST�EM*��V9.1�060 11/�14/2017 A 
  ����CELLSE�T_T  � w$GI_ST�YSEL_P �7T  
7ISO:iRibDiTRA�R|��I_INI; �����bU9A�RTaRSRPNSS1Q23U4567y8Q
TROBQ?ACKSNO� �)�7�E� S�a�o�z�2 3 4 5* 6 7 8aw.n&GINm'D�&� �)%��)4%��)P%���)l%SN�{(O�U��!7� OPT�NA�73�73.:BP<;}a6.:C<;CK;�CaI_DECS�NA�3R�3�TR�Y1��4��4�PTHCN�8D�D>�INCYC@HG��KD�TASKOK�{D�{D�7:�E �U:�Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbH<aRBGSOLA�6�VbG�S�MAx��Vp��Tb@SEGq��T��T�@REQ �d�drG�:Mf�G�JO_HFAUL��Xd�dvgALE@� �g�c�g�cvgE� x�H�dvgNDBR�H<�dgRGAB�Xt�b l�CLM�LIy@   $TYPES�INDEXS�$�$CLASS  ����lq�����apVERSI�ONix ? ���$'61j�r���p��q̛t+ UP0 �x�Style �Select 	�  ��r�uReq. /Echo���yAck�s��sInitiat(�p�r�s�t@�O��a�p���	��  U�����������q�������q���sOption? bit A��p��B����C�Dewcis�cod;���zTryout �mL��Path �segJ�ntin5.�II�yc:��Task OK���!�Manual _opt.r�pA�ԖBޟԖC�� d�ecsn ِ�R�obot int�erlo�"�>� Oisol3��C���i/�"�z�ment���z�ِ����_�s�tatus�	M�H Fault:<��ߧAler���%��p@r 1�z �L��[�m�+�; L�E_COMNT �?�y�    ��䆳�Ŀֿ���� �0�B�T�g�xϊϜ� ������������,� >�P�b�t߆ߘߪ߼�@�����������U�������   ��E�NAB  �� �u�����������MENU>�y��NAME ?%���(%STORE_BOX7FR����F�  %UP�DAT8�>�P�	S�CAN_SLOTk�O�FXp9��N�
CHE0������LABEL��P��SAFEZ **N�$*L6>P bt������ �(:s^� ������/ / 9/$/]/H/Z/l/~/�/ �/�/�/�/�/?? ? 2?D?}?h?�?�?�?�? �?�?�?�?