��   �=�A��*SYST�EM*��V9.1�060 11/�14/2017 A   ����EIP_CF�G_T   �� $VENDO�R  $DE�VTYPE>PR�DCODIREV�ISION>FA�ST_UDP �5 KEEP_IO�_AnSCNpO�PT` Sp $L�OADED� �C�C� IG�ED_wMOD�NET��EXPLCIT_�MS�$HIG�H_SPEE�$EN8021p�DSCP� Hp ��� SPARE��4&ONN.� | $HOS�� !B SC9E�NABL$S�TATN _SZ��S^TOAPI�OTrIgA��R]V�BW&M�oSC.�  7�CXQ�[XX_���CX_��[ kRs�)%'FLA�MU�L�TR�� C_�O�["TOD&IC$i �AS�Z 'sEC{#�#TIMV�CN� Z�&PAT�  @$IDA_FORMA���!�&� �"9"FIG�^�"2�+�!�$ANALOGI� o  4OU� f8FM�$Q�(�4�$$CLA�SS  ����e1��.��.Z0V�ER_c7  ���$'�0 �8. d����� ���0��&p��0���7/ ��ܔ4( 2�;@ �p!192.1�68.1��2  _ 9�k������d!Dummy?  ion1�?����1�1_D gD�:!�l1#��O/BC�onnect<@2HO�O�OvI(�O���J3 _1_C_vKc_���I4q_�_�_V_�_z_<@5�_o#o�_Go�_<@6Qo�o�o6o�oZo<@7�o�o�o'�o<@81as�:<@9������<@A�A�S��w��<@B����Ïf�珊�<@C�!�3�֏W���<@Da�����F�ǟj�<@Eџ����7�ڟ<@FA�q���&���J�<@G���󯖯���<@H!�Q�c����*�<@I����ӿv�����<@J�1�C��g�
�<@Kqϡϳ�V���z�<@L���#���G���<@MQ߁ߓ�6߷�Z�<@�0���ߖߨ�)���nO1�a�s���:�<@P����������<@Q�A�S���w��<@R������f�����<@�a0#����Y��nTa��F�j<@U��7�<@VAq�&�J<@�W����/��A3_K/]/ /�/$/ 6!�_�/�/p/�/�/6! �_+?=?�/a??6!oo �?�?P?�?t?6!�oO O�?AO�?6!O{O�O 0O�OTOfA��O�O�O!_�Of@401_\_n__�_5_GP1�_�_�_�_o�_GP2o<oNo �_rooGP:/�o�o`o �o�oFQ�/-�oQ �oFQ?��@�d FQ�?���1��FQ �?k�}� ���D�FQjO ۏ폐����FQ�OK� ]� ���$�f@5J_�� ͟p�񟔟���_+�=� ��a����*o����P� ѯt����o����A� 䯦�
{���0���T� ��z�����!�Ŀ�� �[�m�ϑ�4Ϧ�Z� ���π�ߤϦ�ʏ;� M���q�ߦ�:��߽�`��߄�f@6���-� ��Q��������@� ��d�ኯ�����1� �����k�}� ���D���j��������$E�IP_SC 2����?. @������ K��f��@ �4F$,ec,kj�� ]�����,> Pbt����� ��//(/:/L/^/6�� � 0�s. �/�/�/>P?t� ,,00?B?T?�� �?�?�?�?�?�?�?O O,O>OPObOtO�O�O��O�O�O�O�O_w!� �/�/?_Q_c_u_�/�/ ??�_�_�_f?x?)o ;oMo_oqo�o�o�o�o �o�o�o%7I [m��:_�� ����_�S��&m&k | �p�����ooʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D��h�W� ������#�5�G�Y�
� �.�����I�v����� ����п�����*� <�N�`�rτϖϨϺ� ����u����&�8�J� ��ϯ��߶���;� ��_��"�4�F�X�j� |������������ ��0�B�T�f�x�� ������������i�{� ����Pbt���ߪ ����(: L^p����� �� //$/��H/7/ l/~/�/'9�/ �/?��)?V?h?z? �?�?�?�?�?�?�?
O O.O@OROdOvO�O�O �O�OU/�O�O__*_ �/�/�/�/�_�_�_? �_??�_oo&o8oJo \ono�o�o�o�o�o�o �o�o"4FX�O |k����I_[_ m_�0�B�T��_�_�� ������ҏ����� ,�>�P�b�t������� ��Ο�����(�� L�^�p�����ʯ ܯ�a�s�	�6�H�Z� l�~�������ƿؿ� ��� �2�D�V�h�z� �Ϟ�5��ϱ�����
� }�������d�v߈��� �����������*� <�N�`�r����� ��������&�8��� \�K���������)�;� M߼�"4�߹�j |������� 0BTfx� �����{�/� ,/>/P/���������/ �/�/AS�/?(?:? L?^?p?�?�?�?�?�? �?�? OO$O6OHOZO lO~O/�O�O�O�O�O ]/o/�/�/D_V_h_�/ �_�/�_�_�_�_�_
o o.o@oRodovo�o�o �o�o�o�o�o�O <+`r��	__ -_�����_�_J� \�n���������ȏڏ ����"�4�F�X�j� |�������ğ[�ן ��0������� ����!�3�ɯ���� ,�>�P�b�t������� ��ο����(�:� L�^�����qϦϸ��� =�O�a�s�$�6�H߻� l�߯�ߢߴ������� ��� �2�D�V�h�z� ������������� ��@�R�d�v����� �|�������g�y�* <N`r���� ���&8J \n���;��� ��/��������j/ |/�/�/�/�/�/ ??0?B?T?f?x?�? �?�?�?�?�?�?OO ,O>O�bOQO�O�O�O ///A/S/__(_�/ L_�/p_�_�_�_�_�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�ooO �o�o 2DV�O�O �O\���G_Y_
� �.�@�R�d�v����� ����Џ����*� <�N�`�r������� ̟ޟ�cu��J� \�n�������ȯگ ����"�4�F�X�j� |�������Ŀֿ��� �ϵ�B�1�f�xϊ� ���!�3������{� ,ߟ�P�b�t߆ߘߪ� ����������(�:� L�^�p�����O� ���� ��$�6��ϻ� ��<�������'�9��� �� 2DVhz �������
 .@Rd��w ���C�U�g�y�*/ </N/����i/�/�/�/ �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?�"OOFOXOjO ��//�O�O�O[/ _/0_B_T_f_x_�_ �_�_�_�_�_�_oo ,o>oPoboto�o�o/O �o�o�o�o�O�O �Op��__� �� ��$�6�H�Z� l�~�������Ə؏� ��� �2�D��oh�W� ������#5GY
� �.���I�v����� ����Я�����*� <�N�`�r��������� ̿޿u���&�8�J� ��ϟ��϶���;� ��_��"�4�F�X�j� |ߎߠ߲��������� ��0�B�T�f�x�� �����������i�{� ����P�b�t����Ϫ� ��������(: L^p����� �� $��H7 l~���'�9�� �/����)/V/h/z/ �/�/�/�/�/�/�/
? ?.?@?R?d?v?�?�? �?�?U�?�?OO*O �����O�O�O/ �O?/�O__&_8_J_ \_n_�_�_�_�_�_�_ �_�_o"o4oFoXo�? |oko�o�o�o�oIO[O mO�o0BT�O�O� �������� ,�>�P�b�t������� ��Ώ�����o(�� L�^�p��o�oʟ ܟ�as	�6�H�Z� l�~�������Ưد� ��� �2�D�V�h�z� ����5�¿�����
� }�������d�vψ��� �����������*� <�N�`�r߄ߖߨߺ� ��������&�8�Ͽ \�K�����)�;� Mϼ��"�4��Ϲ�j� |��������������� 0BTfx� �����{�� ,>P�������� ��A�S��/(/:/ L/^/p/�/�/�/�/�/ �/�/ ??$?6?H?Z? l?~?�?�?�?�?�? ]o��DOVOhO� �O��O�O�O�O�O
_ _._@_R_d_v_�_�_ �_�_�_�_�_oo�? <o+o`oro�o�o	OO -O�o�o�O�OJ \n������ ���"�4�F�X�j� |�������ď[o�׏ ��0��o�o�o�o�� ����!3ɟ���� ,�>�P�b�t������� ��ί����(�:� L�^�����q�����ʿ =�O�a�s�$�6�Hϻ� l�ߟ�Ϣϴ������� ��� �2�D�V�h�z� �ߞ߰��������ߏ� ��@�R�d�v���� �|�������g�y�*� <�N�`�r��������� ������&8J \n���;��� �������j |������� //0/B/T/f/x/�/ �/�/�/�/�/�/?? ,?>?�b?Q?�?�?�? /ASOO(O� LO�pO�O�O�O�O�O �O�O __$_6_H_Z_ l_~_�_�_�_�_�_o? �_�_ o2oDoVo�?�? �?\o�o�o�oGOYO
 .@Rdv�� �������*� <�N�`�r���o���� ̏ޏ��couo�o�oJ� \�n��o�o����ȟڟ ����"�4�F�X�j� |�������į֯��� ����B�1�f�x��� ���!�3�����{� ,ϟ�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸�O� ���� ��$�6奔�� Ϳ<����'�9��� ��� �2�D�V�h�z� ��������������
 .@Rd�߈w ���C�U�g�y�* <N����i��� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/�"??F?X?j? ���?�?�?[ O0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_/? �_�_�_�_oo�?�? �?opo�o�oOO�o �o�o $6HZ l~������ �� �2�D��_h�W� ������#o5oGoYo
� �.��o�oI�v����� ����П�����*� <�N�`�r��������� ̯ޯu���&�8�J� ��Ϗ�󏤿��ȿ;� �_��"�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�x�� �ߋ���������i�{� ����P�b�t������ ����������(�:� L�^�p����������� ���� $��H7 l~���'�9�� ����)Vhz �������
/ /./@/R/d/v/�/�/ �/�/U�/�/??*? �����?�?�? �??�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_�/ |_k_�_�_�_�_I?[? m?�_0oBoTo�?�?�o �o�o�o�o�o�o ,>Pbt��� ������_(�� L�^�p��_�_ooʏ ܏�aoso	�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ����5�¯�����
� }�������d�v����� ���п�����*� <�N�`�rτϖϨϺ� ��������&�8�ϯ \�K߀ߒߤ߶�)�;� M����"�4刺��j� |������������ ��0�B�T�f�x��� ����������{��� ,>P�������ߪ ��A�S��(: L^p����� �� //$/6/H/Z/ l/~/�/�/�/�/�/ ]o��D?V?h?� �?��?�?�?�?�?
O O.O@OROdOvO�O�O �O�O�O�O�O__�/ <_+_`_r_�_�_	?? -?�_�_oo�?�?Jo \ono�o�o�o�o�o�o �o�o"4FXj |����[_�� ��