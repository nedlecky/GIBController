��   v{�A��*SYST�EM*��V9.1�060 11/�14/2017 A   ����UI_CON�FIG_T  �\ J$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�71�ODE�
2�CFOCA �3VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML5C�_wNAM�#DIMC4|:1]ABRIGH83�s oDJ7CH91&U�STO_@  �t @AR$@P�IDD�BC�D*P�AG� ?hAEV�ICE�ISCREVuEF���GN��@$FLAG�@�4&�1  h� 	$PWD_A�CCES� MA�8��LS:1�%)$�LABE� $	Tz j,P�3zR�}	SUSRVI >1  < `oRp*oR�pQPRI��m� t1�PTRI�P�"m�$$CL�A7P �����Q��R��R�P\ S�I��W ? ���$'2 ��,�X�R	_ ,��?2���Ea`NbId�Da����?`�  Gd�o��
 ���Q�o�o�o�o�o	 �o@R dv��)��� ����<�N�`�r� ������7�̏ޏ��� �&���J�\�n����� ��3�ȟڟ����"� 4�ßX�j�|������� A�֯�����0��� T�f�x���������E`TPTX���P����E` s�˸��$/sof�tpart/ge�nlink?he�lp=/md/t�pmenu.dg ¿\�nπϒ�K����� ������ߟ�4�F�X� j�|ߎ�ߟ������� �����B�T�f�x�X�������Q�`p��gbyb�� ($6���������>�ri  �QHad�fcs�fc$d�b�2��k
����dlaha��  ���.�	,�������̷���`���`  ���, +pS ��/#.�F-��c�B 1hR� \��_��� REG V�ED#���wh�olemod.h�tm�	singl��doub��trip�browsF� EWi3��������w��dev.s�lK/�c 1N,	tz/c/� '/�/�/�/�/?#?5?8G?Y?�?� �P�? �?�?�?�?�?OO*O<OFF @�?kO}OLO �O�O�O�F�	}?w?�O __/_A_S_e_w_�_ �_�_�_�_�_�_oo +o=o'UoOo}o�o�o �o�o�o�o�o1 CUgy���� �?�� �2�D�V�h� z������Oԏ���� 
���O�O�d�_�q� ��������˟���� �<�7�I�[������ _o����ٯ����!� 3�E�W�i�{������� ÿտ������X� j�|ώϠϲ������� �����0����f�x� /�A�'��߻������ ��'�P�K�]�o�� ���������ﻯ� �5�G�Y�k�}����� ����������1 CUgyGϴ�� �� 2DVQ� z�[m���ߝ� �//)/;/d/_/q/ �/�/�/�/�/�/�/? ?<?7?I?�i?c?�? �?�?�?�?�?�?O!O 3OEOWOiO{O�O�O�O �O�O�_"_4_F_X_ j_|_�_�_�_��_�_�_�_o0o>j�$U�I_TOPMEN�U 1	`_a�R 
d�aa�A)*def�ault�O�M�*level0 =*�K	 �o�0��oyo�o�btpi�o[23]w8tpst[1x�o5��o�o�or=h58�e01_l.pn�g�y6menu15�y�p�q13�z�rħz�t4�{�sq�� �B�T�f�x������B 0�ŏ׏��������prim=�qp�age,1422,1&�_�q������� ��˟ݟ���%����:�class,5.�c�u���������B�13������h�0���:�53L�@l�~���������:�8[����%�7϶��[�m�ϑϣϵ��I b`_axo�Ϝm߾uq���5�vty*}$qOmf[0,*�	bПc[164w��5�9xuq�K����x2 ��}-��z��w�{i� +�Ϳ߿�������� � K�$�6�H�Z�l�~�� ��������������A�2CUgy� L�����	�� ֯J\n��A�S�1�����//���:�ainedi���O/a/s/�/�/���config=s�ingle&:�wintpF��/�/�/�??����N?��u�gl[55��q�ߑ?dS�p08h�p076y�?�?�72��O�?!O�KO�z�r�z�r4s�xhO�O�x�ڸO*� __'_9_K_]_���_ �_�_�_�_�_�_|_o@#o5oGoYoko�$;�$�doub�%o?�1}3Z�&dual�i38��,4ro�o�oso9�o�n�o�a�oT fx�_����� ���,�>�P�b�t� +�=�>��ȏڏ��� 	�"�4�F�X�j�|��J9?�����1!��O���se��;�q�#�uf����J�H�rO�Oо��.��6#�u7 [���{�������ÿ ������/�A�п e�wωϛϭϿ��ϰ"�1���/�A� S�^�w߉ߛ߭߿��� `�����+�=�O�a� �b��������n���6���-�?�Q�c��$]�74n�������������C�����	�TPTX[209u<=A524�7�b�B51�8x�k��=P0�2�=A��ۤtv�үҀ@2L	0t11�LE��C:�$tre�eview�#�f3���-}381,26 �o////��S/e/w/ �/�/�/</�/�/�/? ?+?vo���5�o� ���?�?�?�/�?�?O@O)O;OF?X?�2q?�2	��O�O�OTO~��1o?�E؞$_6_H_ �6�O��edit �a�O_�_�_�_��� �{_�C�_-o?oQo  Ro~oɕ�o��oW�o �o�o�o1V�o Oy������ �U��6�H�Z�l�~� ���?��Ə؏���� ��2�D�V�h�z���� ��ԟ���
���� @�R�d�v�����)��� Я�������*�N� `�r�������7�̿޿ ���&ϵ�J�\�n� �ϒϤ�Soeo�ωo�� e�!�3�E�W�j�{� �ߟ�߫�������� �/�A�S������ ��������A��,�>� P�b�t���������� ������(:L^ p������  �$6HZl~ ������/ �2/D/V/h/z/�// �/�/�/�/�/
?���� @?��d?��i�?�?�? �?�?�?�?Os?O;O MO_OrO�O�O�O�O{� �O__&_8_J_\_�/ �_�_�_�_�_�_i_�_ o"o4oFoXo�_|o�o �o�o�o�o�owo 0BTf�o��� ���s��,�>� P�b�t��������Ώ ��򏁏�(�:�L�^� p�?1?��U?ʟ1O�O ����#�5�G�Z�k� ٟw�����ůׯ��� ���OV�h�z����� ����¿���
��.� @�Ͽd�vψϚϬϾ� M�������*�<��� N�r߄ߖߨߺ���[� ����&�8�J���n� �������W����� �"�4�F�X���|����������������*default�����*level�8=���5�Se�� �tpst[1�]a	�y�tpio[23����u�@fm�enu7_l.pkng:13?BL5T9g74{u6?L����� 	//f�?/Q/c/u/�/ �/(/�/�/�/�/??�)?�"prim=�:page,74,1.?e?w?�?�?�?��"B6class,13�?�?�?OO0O�?�256OlO~O�O�O�O�#�<ZO�O _`_$_6_9?K218R?�s_�_�_�_�_�O�26��_�_	oo-o?o��$UI_USERVIEW 1�����R 
��Fo��zo�om�o�o�o�o	 �o?Qcu�*� �����o ��$� �_�q�������J�ˏ ݏ���%�ȏI�[� m����<�����4� ���!�3�E��i�{� ������T�կ������ȟ*zoom�0�ZOOMIN ɟ/�ͯ������̿޿ ����&�8�J��n���ϒϤ϶�*ma�xresJ�MAXRESa���e�.�@� R�d�v�ߚ߬߾��� �߅���*�<�N��� _�m���ߧ������� ����8�J�\�n��� #��������������� ��Xj|�� C����� BTfx�5�� �-�//,/>/� b/t/�/�/�/M/�/�/ �/??�'?5?G?�/ o?�?�?�?�?�?? O O$O6OHO�?lO~O�O �O�O_?�O�O�OWO _ 2_D_V_h__�_�_�_ �_�_�_�_
oo.o@o Ro�Q