��   �A��*SYST�EM*��V9.1�060 11/�14/2017 A   ����FSAC_L�ST_T   �8 $CLNT�_NAME �!$IP_ADD�RESSB $A�CCN _LVL  $APPP � 4�$8 A~O  ���z�����o VER�SIONw�  ���$'DEF\ w { ��� ���ENOABLEw ������LIST 1� �  @�!������ 
[.@�d�� ���/�3//W/ */</�/`/�/�/�/�/ �/�/�/??S?&?8? J?�?n?�?�?�?�?�? O�?�?OO"OsOFO�O jO|O�O�O�O�O_�O �O7__\_B_�_f_x_ �_�_�_�W