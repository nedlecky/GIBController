��   ���A��*SYST�EM*��V9.1�060 11/�14/2017 A   ����DCSS_C�PC_T  �$ $COMM�ENT $�ENABLE � $MODJG�RP_NUMKL�\  $U�FRM\] _VT�X M �   �$Y�Z1K �$Z2�STOP�_TYPKDSB�IO�IDXKE�NBL_CALM�D�USE_PR�EDIC? �EL�AY_TIMJS�PEED_CTR�LKOVR_LI�M? p D� L�0��UTOOiL &S>. � 8J\TC�u
!����O�� ZY0  �� �CHG_S{IZ$AP!��E�DIS�M$!�CO+k#c%?#)J�p 	M$JT#�  �&c"�"k#�)�$�'��_SEEXPA�N#N  $SwTAT/ D�FP_BASE �$� K4!Y� 6_V'>H'3��&J- � �m\AXS\UP�LW�7��p�� S5b �,  g?y?�?��?�?���/�'ELEM/� T �B2N�O�GM@CN$SH�A�D6#� $DA�TA)�&e0 �  PJ�@ 2� 
&P5 ɘ� 1U*n   OVSYSoARRZ0ZR)(qViT(�RSkT_ROBOT�X�S�1Ro�U�V$CU�R_��R�$SET�U$"	�0$T P�_MGN�INP_ASSU#�P2! � PCYH�7'` e�f�Hc1�CONFI�G_CHKPE_P�O* mdSHRSTb{gMN#d&T1b�
 RH<H�d� 0 � ld<�KeAVRCFYXHt�5�1� ��W�OA$RܠZSPH/ (7%Q�Q�Q�3�gBOX/ 8�@6!�6!�7 |r�#As�eUIRY@ � ,�FNpE}R@2 $�po �q_S�r��eUIZN/O 0 IF@L*p,�Z_�0�_�08�gu0  @�Q�i�v	�6~�$$�CL`  �S������Q��Q��VERSION���  �w��$' 2 ǈQ   ��p����Ҁ�  ������PC�  �ï���7��W � �Y�I���Da�  �������΢�  d����Cz  ���������� ��W�7��L�I�o� ��������ǟٟ��� �!�3�D�W�h�z��� ����ïկ���
�� /�@�S�d�v�ϛ��� ��ѿ������+�<� O�`�r߄ߗϩϻ�]� ������'���K�9� n��ߥ߷������� ���#�5�F�Y�j�|� �������������� �1�BU�fx���� ����������- >Qbt���� ���/):/M ^/p/�/�����/ � ?/%/[/H?7?l? ~?�/�/�/�/�/�/�? ?!?3?DOW?hOzO�? �?�?�?�?�?�O
_O /O@_SOd_v__�O�O �O�O�_�Oo_+_<o O_`oro�o�_�_�_]o �o�_o'o�oKo9 n��o�o�o�o�o�o �#5F�Yj�|� ���������� �1�B�U�f�x����� ����ӏ�����-� >�Q�b�t��������� ϟͯ���)�:�M� ^�p���������߯ɿ � ��%�[�H�7�l� ~ϑ�����ǿٿ��� �!�3�D�W�h�zߍ� �ϱ���������
�� /�@�S�d�v��߭� ����������+�<� O�`�r�������]� �����'���K�9 n������������� �#5FYj| �������� 1B/Uf/x/�� �����?/-/ >?Q/b?t?�?�/�/�/ �/�?�/O?)?:OM? ^OpO�O�?�?�?�?�O �? _O%O[OH_7_l_ ~_�O�O�O�O�O�O�_ _!_3_DoW_hozo�_ �_�_�_�_�_�o
o /o@Sodv�o�o �o�o��o�+<� O`�r������]��ˏ�r�$DCSS�_CSC 2�#��Q  P�%���D��yd�u�8���\����� ៤���ڟ;���_� "���F���j���ݯ�� �į%��I��m�� B���f�ǿ��뿮�� ҿ�E��i�,ύ�P� ��t����Ϫ����/� ��S��w�:߉߭�p���ߔ��߸���GRPw 2� ���t	��]�H��l�� ������������!� G�2�k�V���z����� ��������
U @yd����� �	�?*cN �r������ ///M/8/q/\/�/ �/�/�/�/�/?�/? 7?"?[?F??�?�?n? �?�?�?�?O�?OEO 0OiO{O�OXO�O�O�O �O�O�O	_/__S_��_GSTAT 2��Y��<� $���  �<�k��Ϲ<�j�?�7���7��7�=���QA�s���dC�j�BP<��U=2T����q4�_�2j�{?�P�Q��P4���Z@в*��۰�q��U�Z��>��|?s��a�)�y?s�zb���m�Y���o�B�D��G
i<dם���R3?rn_�?�P�P��d���(�?r3��>�z?� ����H�D>%��Fk�V`CZa�(��ne�P
�2���+�A�q}��P�D
��
i�=�`�P	��<�^`
�a70G������@�Q �o�_�_�_
i�FX �:��p���y �Y�Q7Y�5[
i
�8� �0�R���f������� ���ҏ��4��d� v������������� �8��L��T�:�L� n�������ү��ʯ� � �"�P�R�����ğ�~�ȿڿ�����꽿�ݷ��]=�h��fq��5��h�w�|6����@e� �D	����]�O-w��z���R��'�d/�R{�>w��Q����G����m=�P}>���"?r��>D��?m�{��B�0��A��B�DA`D�
i���Ծ55?{��e?z��v�c���*>K�?�v�R>8��?�Q��@}r�D�?rh�jH��F]�?z����2
�Q�ҿz��z>>��=�I�v���^��D�"��
i�=�
��{�A<��1�?CоGн�IL~>�6a�?W� N�0�B�T������$� ��(���^�p�
�X� ��l����������� �� �N�4�F���j�|� ����r�x�@���D V0z�������� ����4L jPb����� �t*/<//`/r/L/ �/�/�/�߲���j�|� �Ϡϲ���������� �0�Bߐ�f�x��?�/ �/�/�/|O�O�/�O�O �O�O�O_��6_/ ._l_R_d_�_�_�_�_ �_�_�_ ooo:oho /_�o�O�o�o�o�o (_|oR�oJl �������� � �N�4�V���j� Ə؏������2�D� �<ONO`O??*?<? N?`?r?�?�?�?�?�? �?,OOO��h�z��� &��*�\�6�`�:�L� ����B��ҿ��ʿ� � �"�P�6�Xφ�l� ~ϼϢϴ���ߪ��� F�x�2�|ߎ�h߲��� ���������6�� >�l�R������ ������ ����b�t� N�������������د �������Ɵ؟��� � �2�D�V�h�z�ȯ ����"(��� �������2/D/ ��,�n/@�f/�/�/�/ �/�/�/�/"???X? >?P?r?�?F�L/�?/ �?O*OONO`OV/�? �O�?�O�O�O�O�O_ �O _>_$_6_X_�_l_ �_�_�_HO�_o�_4o Fo ojo|oVot�� >Pbt���� ���d:L ��o�o�o^oP�b��o n���r���Ώ��zO�_ 
��_�@�&�8�Z��� n�����������ڟ� �<��_�~���j��� Ư������P�&�T� �@�n�T�v������� ڿ��ҿ��"��*�X� >�䯚Ϭφ����ϼ� �����"�4��o�o �o"4FXj| ��� ���Z�<� N�`�������0�
�4� � �j�|��dϦ�x� ����������$
, Z@R�v��� ~τ�L�Pb< ��������� 
/�/@/&/X/v/\/ n/�/�/�/�/�/�/� 6?H?"?l?~?X?�?�? �?�����v߈ߚ߬� ����������*�<� N��r���O�?�?�? �?�_�_�?�_�_�_�_ oo� ?Bo?:oxo ^opo�o�o�o�o�o�o �o,$Ft? o ��_����"�4� *o�^��V�x����� ��܏����
�,� Z�@�b���v��ҟ䟀������>�P�^���$DCSS_JP�C 2J�Q ( DGP������������� ��Ư�����c�2� q�V���z�Ͽ���¿ Կ�;�
��q�@�R� dϹψ��Ϭ����%� ��I��*��N�`�r� �ߖ��ߺ����3�� W�&�8�z��n���� ��������A��e� 4���X���|������� ����+��9sB �f����� �9,�P� t����/�� G//(/:/�/^/�/�/ �/�/�/�/?�/ ?B? g?6?H?�?l?~?�?�? �?	O�?-O�?QO OuO DOVO�OzO�O�O�O�O�_��r�S{��L �O___�_��dN_�_ r_�_�_�_�_o�_;o o_o&o�oJo\ono�o �o�o�o%�oI m4�X�|�� �����W��{� B���f�Ï��珮�� ҏ/�����c���P� ��t�џ��������� =��a�(�o�L���p� �������ʯ'��K� �o�6���Z���~�ۿ ����ƿ�5���Y� � }�Dϡ�h��ό��ϰ� ������U��.�@� R߯�v��ߚ��߾�� ��?��c�*��N�`� r��������)��� M��q�8���\����� ������������[ "F�j�����	0TMODE�L 2=[x\��
 <�c
_  �� �q������ �/N/%/7/�/[/m/ /�/�/�/?�/�/8? ?!?3?E?W?i?�O�? c�?�?O�?�?FOO /OAO�OeOwO�O�O�O �O�O�O�OB__+_x_ O_a_�_�_�_�_�_�_ �_�?�?�?oo�oo oo�o�o�o�o�o�o :#5GYk� �������� �l�C�U���=oOo}� ����w����	��-� z�Q�c����������� ϟ�.���d�;�M� _�q�����⯹�˯� ��ŏ��r��[�m� �������ǿٿ&��� �!�n�E�WϤ�{ύ� �ϱ�����"����X� /�Aߎ�)�;�M�{ߍ� c�����0���f�=� O�a�s�������� �����'�9�K��� o�������������( ������GY�} ������� Z1C�gy�� ��/��D//-/ ?/�/9g/y/�/�/ �/?�/?R?)?;?M? �?q?�?�?�?�?O�? �?ONO%O7O�O[OmO �O�O�O�O�/_�/�O �O\_3_E_�_i_{_�_ �_�_�_o�_�_Foo /oAoSoeowo�o�o�o �o�o�o�o+_ �%_Se���� ����'�9���]� o���������ɏۏ� :��#�p�G�Y�k�}� ����w ��ɟ۟H� �1�~�U�g�y�Ư�� ����ӯ�2�	��-� z�Q�c�������濽� Ͽ�.������� ?�QϾ�9ϧϹ����� ��<��%�r�I�[�m� ߑߣ�������&��� �!�3�E�W��{�� ��uχϵ���4���� /�A�S�e��������� ��������f= O�s����� �P����+= �%�����(/ �/^/5/G/Y/�/}/ �/�/�/�/?�/�/? Z?1?C?�?g?y?�?a s��?�?�?	OOhO ?OQO�OuO�O�O�O�O �O_�O_R_)_;_M_ __q_�_�_�_�_o�_ �_o�?`o�?)o;oo o�o�o�o�o�o�o !3E�i{� ������F���/�|�S�e�w����$�DCSS_PST�AT ����݁Q  �  ��� � (�5��Y� �~� |�ހ�������������݅��ߟ�΄SETU�P 	݉BȄ������B�\�ˇT?1SC 2
5�����Cz���������r�CP R��D�DVo��Ho:� L�^�-�������u�ʿ ܿ��$��5�Z� l�;ϐϢϴσ����� ���� �2�D��h�z� Iߞ߰��ߑ�����
� ��.�@�R�!�v��W� ������������ �E�W���8�����n� ��������/�� SewF��|� ���+=a s�T����� /�'/9/K//o/�/ �/b/�/�/�/�/�/? �/5?G?Y?(�}?�?�? (?�?�?�?�?OO1O  OUOgO6OHO�O�O~O �O�O�O�O_-_?__ c_u_�_V_�_�_�_�_ �_o�_)o;oMooqo �o�odo�o�o�o�o �o7I[*� �r?���r�!� 3��W�i�8������� ��Տ���ȏ�/�A� �e�w�F�X������� ����֟+�=�O�� s�����f���ͯ��� ���9�K�]�,��� ����t�ɿۿ�� #Ϫ��Y�k�:Ϗϡ� �ς����������1� C��g�y�Hߝ߯��� ������	���-�?�Q�  �u��V�h����� ������;�M�_�.� ������v������� %��I[m��� �������! 3i{J�� ����/�//A/ S/"/w/�/X/�/�/�/ �/�/??�/=?O?a? 0?�?�?f?x?�?�?�? OO'O�?KO]OoO> �O�O�O>O�O�O�O�O #_5__Y_k_}_L_�_ �_�_�_�_�_o�_1o Coo$oyo�oZo�o�o �o�o�o	�o?Q c2��h��� ���)��M�_�q� @��������Oݏ�v� Џ%�7��[�m��N� ����ǟ������ޟ 3�E��i�{���\��� ïկ�������A� S�"�4�����j���ѿ 㿲���+���O�a� s�Bϗϩ�x�����������$DCSS_�TCPMAP  �����Q @ ���������/����������	���
�����������ɂ  ���������*����������U��������U���� ��!��U"��#��$��%��U&��'��(��)��U*��+��,��-��U.��/��0��1��U2��3��4��5��U6��7��8��9��U:��;��<��=���>��?��@�UI�RO 2��0�n�Z�l�~�� ������������ � 2�D�V�h�z�������V���R�����! 3EWi{��� ������A ��>w����� ��//+/=/O/a/ s/�/�/�/4�/X�/ ??'?9?K?]?o?�? �?�?�?�?�?�?�?O�#O5O�/YO�UIZ�N 2�	 �0�.ҚO�O�Oć�O �O�O_�O4_F_X_'_ |_�_�_c_�_�_�_�_ oo0o�_TofoxoGo �o�o�o�o�o�o�o ,>Pb%��� y�����(�:� 	�^�p���E�����ʏ ��� ��Տ�H�Z��)�~�����aO�UF�RM R��R�8����
���.�@� �d�v�Q�������Я ⯽����<�N�)� r���_�����̿�� ϡ�&�8��\�n�I� �Ϥ�����ϵ���� ��!�F�X�3�|ߎ�i� ����ۿ���ߙ��0� �T�f�A���w�� ���������>�P� +�t���a��������� ����(9^p K������  �6H#l~Y �������� / 2//V/h/C/�/�/y/ �/�/�/�/
?�/.?@? ?d?v?Q?�?�?�� �?�?�?O*OONO`O ;O�O�OqO�O�O�O�O _�O&_8__I_n_�_ [_�_�_�?�_�_�_o "o�_FoXo3o|o�oio �o�o�o�o�o�o0 BfxS���_ ������>�P� +�a�����s���Ώ�� ��ߏ(�:��^�p� K�������